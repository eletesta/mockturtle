module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 ;
  assign n9 = x2 | x3 ;
  assign n10 = x6 & x7 ;
  assign n11 = ~x5 & n10 ;
  assign n12 = x4 & n11 ;
  assign n13 = ~x1 & n12 ;
  assign n14 = ~n9 & n13 ;
  assign n15 = x4 & x5 ;
  assign n16 = x1 | x3 ;
  assign n17 = ( x2 & ~n15 ) | ( x2 & n16 ) | ( ~n15 & n16 ) ;
  assign n18 = n15 | n17 ;
  assign n19 = ~x0 & n18 ;
  assign n20 = ( ~x0 & n14 ) | ( ~x0 & n19 ) | ( n14 & n19 ) ;
  assign n21 = ~x6 & x7 ;
  assign n22 = x2 & x5 ;
  assign n23 = ( x4 & n21 ) | ( x4 & n22 ) | ( n21 & n22 ) ;
  assign n24 = ~x4 & n23 ;
  assign n25 = x6 & ~x7 ;
  assign n26 = ~x5 & n25 ;
  assign n27 = ( x2 & x4 ) | ( x2 & n26 ) | ( x4 & n26 ) ;
  assign n28 = ~x2 & n27 ;
  assign n29 = ~x3 & n28 ;
  assign n30 = ( ~x3 & n24 ) | ( ~x3 & n29 ) | ( n24 & n29 ) ;
  assign n31 = ( ~x0 & x1 ) | ( ~x0 & n30 ) | ( x1 & n30 ) ;
  assign n32 = ( ~x1 & x3 ) | ( ~x1 & x4 ) | ( x3 & x4 ) ;
  assign n33 = x2 & ~n32 ;
  assign n34 = ( x1 & ~x2 ) | ( x1 & n32 ) | ( ~x2 & n32 ) ;
  assign n35 = ( ~x1 & n33 ) | ( ~x1 & n34 ) | ( n33 & n34 ) ;
  assign n36 = ( x2 & x4 ) | ( x2 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n37 = ( x2 & ~x6 ) | ( x2 & n36 ) | ( ~x6 & n36 ) ;
  assign n38 = x2 & ~n37 ;
  assign n39 = n37 | n38 ;
  assign n40 = ( ~x2 & n38 ) | ( ~x2 & n39 ) | ( n38 & n39 ) ;
  assign n41 = ( x1 & n35 ) | ( x1 & ~n40 ) | ( n35 & ~n40 ) ;
  assign n42 = ~x3 & n41 ;
  assign n43 = ( x3 & n35 ) | ( x3 & n42 ) | ( n35 & n42 ) ;
  assign n44 = x0 | n43 ;
  assign n45 = ( x1 & ~n31 ) | ( x1 & n44 ) | ( ~n31 & n44 ) ;
  assign n46 = x3 | x5 ;
  assign n47 = x3 & x4 ;
  assign n48 = x4 & ~x5 ;
  assign n49 = ( n46 & ~n47 ) | ( n46 & n48 ) | ( ~n47 & n48 ) ;
  assign n50 = x2 & ~n49 ;
  assign n51 = ( x1 & ~n49 ) | ( x1 & n50 ) | ( ~n49 & n50 ) ;
  assign n52 = ( ~x1 & x3 ) | ( ~x1 & x5 ) | ( x3 & x5 ) ;
  assign n53 = ( x4 & x5 ) | ( x4 & ~n52 ) | ( x5 & ~n52 ) ;
  assign n54 = ( ~x3 & x4 ) | ( ~x3 & n52 ) | ( x4 & n52 ) ;
  assign n55 = n53 & ~n54 ;
  assign n56 = ~x3 & x5 ;
  assign n57 = ~x4 & n56 ;
  assign n58 = ~x1 & n57 ;
  assign n59 = ~x2 & n58 ;
  assign n60 = ( x3 & x4 ) | ( x3 & ~n32 ) | ( x4 & ~n32 ) ;
  assign n61 = x2 & n32 ;
  assign n62 = ( x1 & n32 ) | ( x1 & n61 ) | ( n32 & n61 ) ;
  assign n63 = n60 & ~n62 ;
  assign n64 = n59 | n63 ;
  assign n65 = ( ~n51 & n55 ) | ( ~n51 & n64 ) | ( n55 & n64 ) ;
  assign n66 = n51 | n65 ;
  assign n67 = ( x2 & x3 ) | ( x2 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n68 = ( x2 & x4 ) | ( x2 & ~n67 ) | ( x4 & ~n67 ) ;
  assign n69 = ( ~x3 & x5 ) | ( ~x3 & n68 ) | ( x5 & n68 ) ;
  assign n70 = n67 | n69 ;
  assign n71 = ( ~n68 & n69 ) | ( ~n68 & n70 ) | ( n69 & n70 ) ;
  assign n72 = ( ~x1 & x6 ) | ( ~x1 & n71 ) | ( x6 & n71 ) ;
  assign n73 = x5 | x6 ;
  assign n74 = x4 & ~n9 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~x1 & n75 ;
  assign n77 = ( ~n71 & n72 ) | ( ~n71 & n76 ) | ( n72 & n76 ) ;
  assign n78 = ( x2 & x5 ) | ( x2 & x6 ) | ( x5 & x6 ) ;
  assign n79 = ( ~x4 & x6 ) | ( ~x4 & n78 ) | ( x6 & n78 ) ;
  assign n80 = x6 & ~n79 ;
  assign n81 = n79 | n80 ;
  assign n82 = ( ~x6 & n80 ) | ( ~x6 & n81 ) | ( n80 & n81 ) ;
  assign n83 = x1 | x7 ;
  assign n84 = ( x3 & n82 ) | ( x3 & n83 ) | ( n82 & n83 ) ;
  assign n85 = n82 & ~n84 ;
  assign n86 = ( ~x0 & n77 ) | ( ~x0 & n85 ) | ( n77 & n85 ) ;
  assign n87 = ~n66 & n86 ;
  assign n88 = ( ~x0 & n66 ) | ( ~x0 & n87 ) | ( n66 & n87 ) ;
  assign n89 = ( x3 & x5 ) | ( x3 & x6 ) | ( x5 & x6 ) ;
  assign n90 = x3 & n89 ;
  assign n91 = ( x2 & ~x3 ) | ( x2 & n89 ) | ( ~x3 & n89 ) ;
  assign n92 = ~n89 & n91 ;
  assign n93 = n90 | n92 ;
  assign n94 = ~x1 & n93 ;
  assign n95 = x2 | n73 ;
  assign n96 = ( ~x1 & x3 ) | ( ~x1 & n95 ) | ( x3 & n95 ) ;
  assign n97 = x1 | n96 ;
  assign n98 = ( x2 & ~x3 ) | ( x2 & x5 ) | ( ~x3 & x5 ) ;
  assign n99 = ( x2 & x3 ) | ( x2 & ~x6 ) | ( x3 & ~x6 ) ;
  assign n100 = n98 | n99 ;
  assign n101 = ( x3 & ~x5 ) | ( x3 & n100 ) | ( ~x5 & n100 ) ;
  assign n102 = x4 | n101 ;
  assign n103 = ~x2 & x3 ;
  assign n104 = x5 & x6 ;
  assign n105 = n103 & n104 ;
  assign n106 = x4 & ~n105 ;
  assign n107 = n102 & ~n106 ;
  assign n108 = x1 | n107 ;
  assign n109 = x4 | n73 ;
  assign n110 = n103 & ~n109 ;
  assign n111 = x1 & ~n110 ;
  assign n112 = n108 & ~n111 ;
  assign n113 = n97 & ~n112 ;
  assign n114 = ( ~n93 & n94 ) | ( ~n93 & n113 ) | ( n94 & n113 ) ;
  assign n115 = ( x1 & x2 ) | ( x1 & x4 ) | ( x2 & x4 ) ;
  assign n116 = ( x3 & x6 ) | ( x3 & n115 ) | ( x6 & n115 ) ;
  assign n117 = ( x5 & ~x6 ) | ( x5 & n116 ) | ( ~x6 & n116 ) ;
  assign n118 = ( x3 & x5 ) | ( x3 & ~n116 ) | ( x5 & ~n116 ) ;
  assign n119 = n117 & ~n118 ;
  assign n120 = ~x2 & x4 ;
  assign n121 = x3 & n120 ;
  assign n122 = x5 & n21 ;
  assign n123 = n121 & n122 ;
  assign n124 = ( ~x4 & x6 ) | ( ~x4 & x7 ) | ( x6 & x7 ) ;
  assign n125 = ( x2 & ~x6 ) | ( x2 & n124 ) | ( ~x6 & n124 ) ;
  assign n126 = ( ~x4 & x7 ) | ( ~x4 & n125 ) | ( x7 & n125 ) ;
  assign n127 = ~n124 & n126 ;
  assign n128 = ( ~n125 & n126 ) | ( ~n125 & n127 ) | ( n126 & n127 ) ;
  assign n129 = ( x3 & ~x5 ) | ( x3 & n128 ) | ( ~x5 & n128 ) ;
  assign n130 = ( n29 & n128 ) | ( n29 & ~n129 ) | ( n128 & ~n129 ) ;
  assign n131 = x1 & ~n9 ;
  assign n132 = ( ~n15 & n21 ) | ( ~n15 & n131 ) | ( n21 & n131 ) ;
  assign n133 = n15 & n132 ;
  assign n134 = ( ~n123 & n130 ) | ( ~n123 & n133 ) | ( n130 & n133 ) ;
  assign n135 = x1 & ~n133 ;
  assign n136 = ( n123 & n134 ) | ( n123 & ~n135 ) | ( n134 & ~n135 ) ;
  assign n137 = ( ~x0 & n119 ) | ( ~x0 & n136 ) | ( n119 & n136 ) ;
  assign n138 = n114 & n137 ;
  assign n139 = ( x0 & n114 ) | ( x0 & ~n138 ) | ( n114 & ~n138 ) ;
  assign n140 = x3 & x5 ;
  assign n141 = x5 & ~x7 ;
  assign n142 = ( x1 & n140 ) | ( x1 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( ~x1 & x7 ) | ( ~x1 & n142 ) | ( x7 & n142 ) ;
  assign n144 = ( ~x5 & n140 ) | ( ~x5 & n143 ) | ( n140 & n143 ) ;
  assign n145 = ( ~n140 & n142 ) | ( ~n140 & n144 ) | ( n142 & n144 ) ;
  assign n146 = ~x3 & n25 ;
  assign n147 = ( x1 & ~x5 ) | ( x1 & n146 ) | ( ~x5 & n146 ) ;
  assign n148 = ~x1 & n147 ;
  assign n149 = x6 & ~n148 ;
  assign n150 = ( n145 & n148 ) | ( n145 & ~n149 ) | ( n148 & ~n149 ) ;
  assign n151 = x4 & ~n150 ;
  assign n152 = ( x3 & x6 ) | ( x3 & x7 ) | ( x6 & x7 ) ;
  assign n153 = ( ~x3 & x5 ) | ( ~x3 & n152 ) | ( x5 & n152 ) ;
  assign n154 = ( x6 & x7 ) | ( x6 & n153 ) | ( x7 & n153 ) ;
  assign n155 = ~n152 & n154 ;
  assign n156 = ( ~n153 & n154 ) | ( ~n153 & n155 ) | ( n154 & n155 ) ;
  assign n157 = ~x1 & n156 ;
  assign n158 = x4 | n157 ;
  assign n159 = ~n151 & n158 ;
  assign n160 = x2 | n159 ;
  assign n161 = ( x5 & ~x6 ) | ( x5 & x7 ) | ( ~x6 & x7 ) ;
  assign n162 = ~x7 & n161 ;
  assign n163 = ( x4 & ~x5 ) | ( x4 & n162 ) | ( ~x5 & n162 ) ;
  assign n164 = ( n161 & n162 ) | ( n161 & n163 ) | ( n162 & n163 ) ;
  assign n165 = x3 | n164 ;
  assign n166 = ~x4 & n11 ;
  assign n167 = x3 & ~n166 ;
  assign n168 = n165 & ~n167 ;
  assign n169 = ~x1 & n168 ;
  assign n170 = x2 & ~n169 ;
  assign n171 = n160 & ~n170 ;
  assign n172 = ( ~x1 & x2 ) | ( ~x1 & n9 ) | ( x2 & n9 ) ;
  assign n173 = ( x1 & x2 ) | ( x1 & ~n9 ) | ( x2 & ~n9 ) ;
  assign n174 = ( ~x2 & n172 ) | ( ~x2 & n173 ) | ( n172 & n173 ) ;
  assign n175 = ( x5 & x6 ) | ( x5 & n174 ) | ( x6 & n174 ) ;
  assign n176 = ( x4 & ~x6 ) | ( x4 & n175 ) | ( ~x6 & n175 ) ;
  assign n177 = ( x4 & x5 ) | ( x4 & ~n175 ) | ( x5 & ~n175 ) ;
  assign n178 = n176 & ~n177 ;
  assign n179 = ~x1 & x2 ;
  assign n180 = ~x1 & x4 ;
  assign n181 = ( n120 & n179 ) | ( n120 & ~n180 ) | ( n179 & ~n180 ) ;
  assign n182 = ( ~x3 & x6 ) | ( ~x3 & n181 ) | ( x6 & n181 ) ;
  assign n183 = ( x5 & ~x6 ) | ( x5 & n182 ) | ( ~x6 & n182 ) ;
  assign n184 = ( x3 & ~x5 ) | ( x3 & n182 ) | ( ~x5 & n182 ) ;
  assign n185 = n183 & n184 ;
  assign n186 = x1 & ~x2 ;
  assign n187 = x1 | n9 ;
  assign n188 = ( ~x1 & n186 ) | ( ~x1 & n187 ) | ( n186 & n187 ) ;
  assign n189 = ( x4 & ~x6 ) | ( x4 & n188 ) | ( ~x6 & n188 ) ;
  assign n190 = ( ~x5 & x6 ) | ( ~x5 & n189 ) | ( x6 & n189 ) ;
  assign n191 = ( ~x4 & x5 ) | ( ~x4 & n189 ) | ( x5 & n189 ) ;
  assign n192 = n190 | n191 ;
  assign n193 = x4 | x6 ;
  assign n194 = ( ~x2 & x4 ) | ( ~x2 & x6 ) | ( x4 & x6 ) ;
  assign n195 = ( x3 & x4 ) | ( x3 & n194 ) | ( x4 & n194 ) ;
  assign n196 = n194 & n195 ;
  assign n197 = n193 & ~n196 ;
  assign n198 = x1 & ~n197 ;
  assign n199 = x3 & ~x6 ;
  assign n200 = x4 & ~x6 ;
  assign n201 = ( ~x5 & x6 ) | ( ~x5 & n200 ) | ( x6 & n200 ) ;
  assign n202 = ( x3 & ~x5 ) | ( x3 & n200 ) | ( ~x5 & n200 ) ;
  assign n203 = ( n199 & n201 ) | ( n199 & ~n202 ) | ( n201 & ~n202 ) ;
  assign n204 = x2 & n203 ;
  assign n205 = x1 | n204 ;
  assign n206 = ~n198 & n205 ;
  assign n207 = n192 & ~n206 ;
  assign n208 = ( n178 & ~n185 ) | ( n178 & n207 ) | ( ~n185 & n207 ) ;
  assign n209 = ~n178 & n208 ;
  assign n210 = x0 | n209 ;
  assign n211 = ( x0 & ~n171 ) | ( x0 & n210 ) | ( ~n171 & n210 ) ;
  assign n212 = ( ~x0 & x2 ) | ( ~x0 & n16 ) | ( x2 & n16 ) ;
  assign n213 = x0 | n212 ;
  assign n214 = x5 | n213 ;
  assign n215 = ( ~x4 & x6 ) | ( ~x4 & n214 ) | ( x6 & n214 ) ;
  assign n216 = x4 | n215 ;
  assign n217 = x7 | n216 ;
  assign n218 = x5 & ~x6 ;
  assign n219 = ~x7 & n218 ;
  assign n220 = x5 | n219 ;
  assign n221 = x3 | x4 ;
  assign n222 = ( ~n219 & n220 ) | ( ~n219 & n221 ) | ( n220 & n221 ) ;
  assign n223 = x1 | n222 ;
  assign n224 = ( ~x0 & x2 ) | ( ~x0 & n223 ) | ( x2 & n223 ) ;
  assign n225 = x0 | n224 ;
  assign n226 = ( x4 & ~x5 ) | ( x4 & x6 ) | ( ~x5 & x6 ) ;
  assign n227 = ( ~x4 & x5 ) | ( ~x4 & n226 ) | ( x5 & n226 ) ;
  assign n228 = x7 & ~n226 ;
  assign n229 = ( x6 & ~n226 ) | ( x6 & n228 ) | ( ~n226 & n228 ) ;
  assign n230 = n227 & ~n229 ;
  assign n231 = ( x2 & n16 ) | ( x2 & ~n230 ) | ( n16 & ~n230 ) ;
  assign n232 = n230 | n231 ;
  assign n233 = x0 | n232 ;
  assign n234 = ( x3 & x5 ) | ( x3 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n235 = ( x3 & x4 ) | ( x3 & ~n234 ) | ( x4 & ~n234 ) ;
  assign n236 = ( ~x5 & x7 ) | ( ~x5 & n235 ) | ( x7 & n235 ) ;
  assign n237 = n234 | n236 ;
  assign n238 = ( ~n235 & n236 ) | ( ~n235 & n237 ) | ( n236 & n237 ) ;
  assign n239 = x6 & ~n238 ;
  assign n240 = n26 & ~n221 ;
  assign n241 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n242 = x3 & ~n241 ;
  assign n243 = ( x6 & n56 ) | ( x6 & n242 ) | ( n56 & n242 ) ;
  assign n244 = n242 | n243 ;
  assign n245 = n240 | n244 ;
  assign n246 = ( n238 & n239 ) | ( n238 & ~n245 ) | ( n239 & ~n245 ) ;
  assign n247 = x0 | x2 ;
  assign n248 = ( x1 & ~n246 ) | ( x1 & n247 ) | ( ~n246 & n247 ) ;
  assign n249 = n246 | n248 ;
  assign n250 = ~x5 & x6 ;
  assign n251 = x6 & ~n250 ;
  assign n252 = x4 & n251 ;
  assign n253 = ( x3 & n250 ) | ( x3 & ~n251 ) | ( n250 & ~n251 ) ;
  assign n254 = ( x5 & ~n252 ) | ( x5 & n253 ) | ( ~n252 & n253 ) ;
  assign n255 = ( x3 & ~x5 ) | ( x3 & x6 ) | ( ~x5 & x6 ) ;
  assign n256 = ( x3 & ~x7 ) | ( x3 & n255 ) | ( ~x7 & n255 ) ;
  assign n257 = x3 & ~n256 ;
  assign n258 = n256 | n257 ;
  assign n259 = ( ~x3 & n257 ) | ( ~x3 & n258 ) | ( n257 & n258 ) ;
  assign n260 = x4 & ~n259 ;
  assign n261 = ( x5 & x6 ) | ( x5 & x7 ) | ( x6 & x7 ) ;
  assign n262 = ~x6 & n261 ;
  assign n263 = ( ~x5 & n261 ) | ( ~x5 & n262 ) | ( n261 & n262 ) ;
  assign n264 = ~x3 & n263 ;
  assign n265 = x4 | n264 ;
  assign n266 = ~n260 & n265 ;
  assign n267 = x2 & ~x3 ;
  assign n268 = ~x4 & x5 ;
  assign n269 = ( x3 & x4 ) | ( x3 & n268 ) | ( x4 & n268 ) ;
  assign n270 = ( ~x2 & x3 ) | ( ~x2 & n269 ) | ( x3 & n269 ) ;
  assign n271 = ( n267 & ~n269 ) | ( n267 & n270 ) | ( ~n269 & n270 ) ;
  assign n272 = ( n254 & n266 ) | ( n254 & n271 ) | ( n266 & n271 ) ;
  assign n273 = x2 & ~n271 ;
  assign n274 = ( n254 & ~n272 ) | ( n254 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = x1 | n274 ;
  assign n276 = x0 | n275 ;
  assign n277 = ( x3 & ~x4 ) | ( x3 & x6 ) | ( ~x4 & x6 ) ;
  assign n278 = ( x3 & ~x7 ) | ( x3 & n277 ) | ( ~x7 & n277 ) ;
  assign n279 = x3 & ~n278 ;
  assign n280 = n278 | n279 ;
  assign n281 = ( ~x3 & n279 ) | ( ~x3 & n280 ) | ( n279 & n280 ) ;
  assign n282 = x5 & ~n281 ;
  assign n283 = ( x4 & x7 ) | ( x4 & n200 ) | ( x7 & n200 ) ;
  assign n284 = ( ~x4 & x7 ) | ( ~x4 & n200 ) | ( x7 & n200 ) ;
  assign n285 = ( x4 & ~n283 ) | ( x4 & n284 ) | ( ~n283 & n284 ) ;
  assign n286 = x3 | n285 ;
  assign n287 = ~x5 & n286 ;
  assign n288 = n282 | n287 ;
  assign n289 = ~x2 & n288 ;
  assign n290 = n219 & ~n221 ;
  assign n291 = x2 & ~n290 ;
  assign n292 = n289 | n291 ;
  assign n293 = ( x0 & x1 ) | ( x0 & ~n292 ) | ( x1 & ~n292 ) ;
  assign n294 = ( x1 & ~x3 ) | ( x1 & x5 ) | ( ~x3 & x5 ) ;
  assign n295 = ( x2 & ~x5 ) | ( x2 & n294 ) | ( ~x5 & n294 ) ;
  assign n296 = ( ~x1 & x5 ) | ( ~x1 & n295 ) | ( x5 & n295 ) ;
  assign n297 = ~n294 & n296 ;
  assign n298 = x2 & ~n297 ;
  assign n299 = ( n295 & n297 ) | ( n295 & ~n298 ) | ( n297 & ~n298 ) ;
  assign n300 = x4 & n299 ;
  assign n301 = x2 & x4 ;
  assign n302 = ( x1 & x3 ) | ( x1 & n301 ) | ( x3 & n301 ) ;
  assign n303 = ~x1 & n302 ;
  assign n304 = x4 & x6 ;
  assign n305 = x1 & ~x6 ;
  assign n306 = x1 & n221 ;
  assign n307 = ( n304 & n305 ) | ( n304 & ~n306 ) | ( n305 & ~n306 ) ;
  assign n308 = x5 & n307 ;
  assign n309 = ~x2 & n308 ;
  assign n310 = n303 | n309 ;
  assign n311 = ( n299 & ~n300 ) | ( n299 & n310 ) | ( ~n300 & n310 ) ;
  assign n312 = ~x0 & n311 ;
  assign n313 = ( n292 & n293 ) | ( n292 & ~n312 ) | ( n293 & ~n312 ) ;
  assign n314 = ( x1 & x5 ) | ( x1 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n315 = ( x1 & x4 ) | ( x1 & ~n250 ) | ( x4 & ~n250 ) ;
  assign n316 = ~n314 & n315 ;
  assign n317 = ( ~x2 & x3 ) | ( ~x2 & n316 ) | ( x3 & n316 ) ;
  assign n318 = ( ~x5 & n180 ) | ( ~x5 & n304 ) | ( n180 & n304 ) ;
  assign n319 = ( x5 & x6 ) | ( x5 & ~n180 ) | ( x6 & ~n180 ) ;
  assign n320 = ( ~x6 & n318 ) | ( ~x6 & n319 ) | ( n318 & n319 ) ;
  assign n321 = ( x2 & x3 ) | ( x2 & ~n320 ) | ( x3 & ~n320 ) ;
  assign n322 = n317 & ~n321 ;
  assign n323 = x1 | x2 ;
  assign n324 = x2 & ~n16 ;
  assign n325 = ( ~x2 & n323 ) | ( ~x2 & n324 ) | ( n323 & n324 ) ;
  assign n326 = ( x4 & x6 ) | ( x4 & n325 ) | ( x6 & n325 ) ;
  assign n327 = ( x5 & ~x6 ) | ( x5 & n326 ) | ( ~x6 & n326 ) ;
  assign n328 = ( x4 & x5 ) | ( x4 & ~n326 ) | ( x5 & ~n326 ) ;
  assign n329 = n327 & ~n328 ;
  assign n330 = ( x4 & x5 ) | ( x4 & ~n294 ) | ( x5 & ~n294 ) ;
  assign n331 = ( ~x1 & x3 ) | ( ~x1 & n330 ) | ( x3 & n330 ) ;
  assign n332 = n294 | n331 ;
  assign n333 = ( ~n330 & n331 ) | ( ~n330 & n332 ) | ( n331 & n332 ) ;
  assign n334 = ~x2 & n333 ;
  assign n335 = x3 & ~x4 ;
  assign n336 = ~x1 & n335 ;
  assign n337 = x2 & ~n336 ;
  assign n338 = n334 | n337 ;
  assign n339 = ~n329 & n338 ;
  assign n340 = ~n322 & n339 ;
  assign n341 = ( x1 & x3 ) | ( x1 & ~x7 ) | ( x3 & ~x7 ) ;
  assign n342 = ( x1 & x6 ) | ( x1 & ~n341 ) | ( x6 & ~n341 ) ;
  assign n343 = ( ~x3 & x7 ) | ( ~x3 & n342 ) | ( x7 & n342 ) ;
  assign n344 = n341 | n343 ;
  assign n345 = ( ~n342 & n343 ) | ( ~n342 & n344 ) | ( n343 & n344 ) ;
  assign n346 = x4 & ~n345 ;
  assign n347 = ( ~x3 & x6 ) | ( ~x3 & x7 ) | ( x6 & x7 ) ;
  assign n348 = ( x4 & x6 ) | ( x4 & x7 ) | ( x6 & x7 ) ;
  assign n349 = n347 & ~n348 ;
  assign n350 = n346 | n349 ;
  assign n351 = ( ~x1 & n346 ) | ( ~x1 & n350 ) | ( n346 & n350 ) ;
  assign n352 = ( x2 & ~x5 ) | ( x2 & n351 ) | ( ~x5 & n351 ) ;
  assign n353 = ~x5 & n335 ;
  assign n354 = ( x1 & n21 ) | ( x1 & n353 ) | ( n21 & n353 ) ;
  assign n355 = ~x1 & n354 ;
  assign n356 = ~x2 & n355 ;
  assign n357 = ( n351 & ~n352 ) | ( n351 & n356 ) | ( ~n352 & n356 ) ;
  assign n358 = ~x3 & x4 ;
  assign n359 = ( x5 & ~x7 ) | ( x5 & n358 ) | ( ~x7 & n358 ) ;
  assign n360 = ( x4 & x5 ) | ( x4 & ~n358 ) | ( x5 & ~n358 ) ;
  assign n361 = ( x3 & x7 ) | ( x3 & ~n360 ) | ( x7 & ~n360 ) ;
  assign n362 = n359 | n361 ;
  assign n363 = ( ~x6 & n179 ) | ( ~x6 & n362 ) | ( n179 & n362 ) ;
  assign n364 = ~n362 & n363 ;
  assign n365 = ( ~x0 & n357 ) | ( ~x0 & n364 ) | ( n357 & n364 ) ;
  assign n366 = n340 & n365 ;
  assign n367 = ( x0 & n340 ) | ( x0 & ~n366 ) | ( n340 & ~n366 ) ;
  assign n368 = ( x2 & ~x4 ) | ( x2 & x7 ) | ( ~x4 & x7 ) ;
  assign n369 = ~x3 & x6 ;
  assign n370 = ( n56 & n250 ) | ( n56 & ~n369 ) | ( n250 & ~n369 ) ;
  assign n371 = x2 | x7 ;
  assign n372 = ( ~x4 & n370 ) | ( ~x4 & n371 ) | ( n370 & n371 ) ;
  assign n373 = ~n368 & n372 ;
  assign n374 = ( x2 & n21 ) | ( x2 & n353 ) | ( n21 & n353 ) ;
  assign n375 = ~x2 & n374 ;
  assign n376 = x6 | x7 ;
  assign n377 = x2 & ~x4 ;
  assign n378 = ~x2 & x5 ;
  assign n379 = x3 & ~n378 ;
  assign n380 = ( n47 & n377 ) | ( n47 & ~n379 ) | ( n377 & ~n379 ) ;
  assign n381 = ( x6 & x7 ) | ( x6 & ~n380 ) | ( x7 & ~n380 ) ;
  assign n382 = ( n375 & n376 ) | ( n375 & ~n381 ) | ( n376 & ~n381 ) ;
  assign n383 = n373 | n382 ;
  assign n384 = x1 | n383 ;
  assign n385 = n10 & n15 ;
  assign n386 = n103 & n385 ;
  assign n387 = x1 & ~n386 ;
  assign n388 = n384 & ~n387 ;
  assign n389 = ( x5 & x6 ) | ( x5 & ~n277 ) | ( x6 & ~n277 ) ;
  assign n390 = ( ~x3 & x5 ) | ( ~x3 & n277 ) | ( x5 & n277 ) ;
  assign n391 = n389 & ~n390 ;
  assign n392 = x2 & ~n391 ;
  assign n393 = x3 | n109 ;
  assign n394 = ~x2 & n393 ;
  assign n395 = n392 | n394 ;
  assign n396 = ~x1 & n395 ;
  assign n397 = ~x4 & n104 ;
  assign n398 = ~n9 & n397 ;
  assign n399 = x1 & ~n398 ;
  assign n400 = n396 | n399 ;
  assign n401 = ( x3 & x7 ) | ( x3 & n15 ) | ( x7 & n15 ) ;
  assign n402 = ( x3 & x7 ) | ( x3 & ~n15 ) | ( x7 & ~n15 ) ;
  assign n403 = ( x4 & x5 ) | ( x4 & n402 ) | ( x5 & n402 ) ;
  assign n404 = ~n401 & n403 ;
  assign n405 = x2 | n404 ;
  assign n406 = ~x5 & x7 ;
  assign n407 = x4 & n406 ;
  assign n408 = x3 & n407 ;
  assign n409 = x2 & ~n408 ;
  assign n410 = n405 & ~n409 ;
  assign n411 = n179 & n353 ;
  assign n412 = ( ~x1 & n410 ) | ( ~x1 & n411 ) | ( n410 & n411 ) ;
  assign n413 = x2 | x4 ;
  assign n414 = ( x2 & ~x3 ) | ( x2 & n413 ) | ( ~x3 & n413 ) ;
  assign n415 = ( x1 & n411 ) | ( x1 & n414 ) | ( n411 & n414 ) ;
  assign n416 = n412 | n415 ;
  assign n417 = ( x0 & n400 ) | ( x0 & ~n416 ) | ( n400 & ~n416 ) ;
  assign n418 = n388 | n417 ;
  assign n419 = ( x0 & ~n388 ) | ( x0 & n418 ) | ( ~n388 & n418 ) ;
  assign y0 = ~x0 ;
  assign y1 = ~x0 ;
  assign y2 = ~x0 ;
  assign y3 = n20 ;
  assign y4 = ~n45 ;
  assign y5 = n88 ;
  assign y6 = ~n139 ;
  assign y7 = ~n211 ;
  assign y8 = ~n217 ;
  assign y9 = ~n225 ;
  assign y10 = ~n233 ;
  assign y11 = ~n249 ;
  assign y12 = ~n276 ;
  assign y13 = ~n313 ;
  assign y14 = ~n367 ;
  assign y15 = ~n419 ;
endmodule
