module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 ;
  assign n7 = ( x1 & x2 ) | ( x1 & x3 ) | ( x2 & x3 ) ;
  assign n8 = x4 & ~n7 ;
  assign n9 = ( x1 & x4 ) | ( x1 & ~n8 ) | ( x4 & ~n8 ) ;
  assign n10 = x0 & n9 ;
  assign n11 = x1 & ~x2 ;
  assign n12 = x3 & ~x4 ;
  assign n13 = ( x2 & ~x3 ) | ( x2 & n12 ) | ( ~x3 & n12 ) ;
  assign n14 = ( ~x1 & x2 ) | ( ~x1 & n13 ) | ( x2 & n13 ) ;
  assign n15 = ( n11 & ~n13 ) | ( n11 & n14 ) | ( ~n13 & n14 ) ;
  assign n16 = x0 & ~n15 ;
  assign n17 = ( x0 & x3 ) | ( x0 & x4 ) | ( x3 & x4 ) ;
  assign n18 = ( x0 & x3 ) | ( x0 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n19 = n17 & ~n18 ;
  assign n20 = x2 & ~x4 ;
  assign n21 = x3 & n20 ;
  assign n22 = x1 | x3 ;
  assign n23 = ( x0 & ~x2 ) | ( x0 & n22 ) | ( ~x2 & n22 ) ;
  assign n24 = ( x0 & x3 ) | ( x0 & ~n22 ) | ( x3 & ~n22 ) ;
  assign n25 = ( x1 & ~n23 ) | ( x1 & n24 ) | ( ~n23 & n24 ) ;
  assign n26 = ( x0 & ~x1 ) | ( x0 & n25 ) | ( ~x1 & n25 ) ;
  assign n27 = n21 & ~n26 ;
  assign n28 = ( n21 & n25 ) | ( n21 & ~n27 ) | ( n25 & ~n27 ) ;
  assign n29 = ( x1 & ~x2 ) | ( x1 & n28 ) | ( ~x2 & n28 ) ;
  assign n30 = n19 & ~n29 ;
  assign n31 = ( n19 & n28 ) | ( n19 & ~n30 ) | ( n28 & ~n30 ) ;
  assign n32 = ( x1 & ~x3 ) | ( x1 & x5 ) | ( ~x3 & x5 ) ;
  assign n33 = ( x2 & ~x5 ) | ( x2 & n32 ) | ( ~x5 & n32 ) ;
  assign n34 = ( x1 & x2 ) | ( x1 & ~n32 ) | ( x2 & ~n32 ) ;
  assign n35 = n33 & ~n34 ;
  assign n36 = x0 & ~n35 ;
  assign n37 = ~x2 & x3 ;
  assign n38 = ~x5 & n37 ;
  assign n39 = x1 & n38 ;
  assign n40 = x0 | n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = ~x4 & n41 ;
  assign n43 = ( x0 & ~x2 ) | ( x0 & x3 ) | ( ~x2 & x3 ) ;
  assign n44 = ( ~x0 & x1 ) | ( ~x0 & n43 ) | ( x1 & n43 ) ;
  assign n45 = ( ~x2 & x3 ) | ( ~x2 & n44 ) | ( x3 & n44 ) ;
  assign n46 = ~n43 & n45 ;
  assign n47 = ( ~n44 & n45 ) | ( ~n44 & n46 ) | ( n45 & n46 ) ;
  assign n48 = ( x1 & ~x2 ) | ( x1 & x3 ) | ( ~x2 & x3 ) ;
  assign n49 = x1 & x4 ;
  assign n50 = ( x3 & ~n48 ) | ( x3 & n49 ) | ( ~n48 & n49 ) ;
  assign n51 = ( ~x4 & n48 ) | ( ~x4 & n50 ) | ( n48 & n50 ) ;
  assign n52 = ( ~x3 & n50 ) | ( ~x3 & n51 ) | ( n50 & n51 ) ;
  assign n53 = x0 & ~n52 ;
  assign n54 = ~x4 & n37 ;
  assign n55 = x1 & n54 ;
  assign n56 = x0 | n55 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = n47 | n57 ;
  assign n59 = ( n41 & ~n42 ) | ( n41 & n58 ) | ( ~n42 & n58 ) ;
  assign n60 = ( x1 & x2 ) | ( x1 & ~x5 ) | ( x2 & ~x5 ) ;
  assign n61 = n7 | n60 ;
  assign n62 = x5 & n61 ;
  assign n63 = ( ~n7 & n61 ) | ( ~n7 & n62 ) | ( n61 & n62 ) ;
  assign n64 = x4 & ~n63 ;
  assign n65 = ~x3 & x5 ;
  assign n66 = ( x1 & x5 ) | ( x1 & n65 ) | ( x5 & n65 ) ;
  assign n67 = x2 & n66 ;
  assign n68 = x4 | n67 ;
  assign n69 = ~n64 & n68 ;
  assign n70 = ~x0 & n69 ;
  assign n71 = x4 & ~x5 ;
  assign n72 = ~x0 & x1 ;
  assign n73 = ~x2 & n72 ;
  assign n74 = x3 & n73 ;
  assign n75 = n71 & n74 ;
  assign n76 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n77 = x2 | n76 ;
  assign n78 = ( x0 & ~x3 ) | ( x0 & n76 ) | ( ~x3 & n76 ) ;
  assign n79 = x2 & n78 ;
  assign n80 = n77 & ~n79 ;
  assign n81 = x4 & ~n80 ;
  assign n82 = x1 | x2 ;
  assign n83 = ( ~x1 & n11 ) | ( ~x1 & n82 ) | ( n11 & n82 ) ;
  assign n84 = x3 & n83 ;
  assign n85 = x4 | n84 ;
  assign n86 = ~n81 & n85 ;
  assign n87 = n75 | n86 ;
  assign n88 = ( n69 & ~n70 ) | ( n69 & n87 ) | ( ~n70 & n87 ) ;
  assign n89 = x2 | x3 ;
  assign n90 = ( x0 & ~x2 ) | ( x0 & n89 ) | ( ~x2 & n89 ) ;
  assign n91 = ( x0 & ~x1 ) | ( x0 & n89 ) | ( ~x1 & n89 ) ;
  assign n92 = ( n11 & ~n90 ) | ( n11 & n91 ) | ( ~n90 & n91 ) ;
  assign n93 = ~x4 & n92 ;
  assign n94 = x2 & ~x3 ;
  assign n95 = ( x0 & ~x4 ) | ( x0 & n94 ) | ( ~x4 & n94 ) ;
  assign n96 = ~x0 & n95 ;
  assign n97 = ( x0 & ~x3 ) | ( x0 & x5 ) | ( ~x3 & x5 ) ;
  assign n98 = ( ~x1 & x5 ) | ( ~x1 & n97 ) | ( x5 & n97 ) ;
  assign n99 = x5 & ~n98 ;
  assign n100 = n98 | n99 ;
  assign n101 = ( ~x5 & n99 ) | ( ~x5 & n100 ) | ( n99 & n100 ) ;
  assign n102 = ~x2 & n101 ;
  assign n103 = ~x2 & x5 ;
  assign n104 = ( x0 & x1 ) | ( x0 & n103 ) | ( x1 & n103 ) ;
  assign n105 = ~x1 & n104 ;
  assign n106 = ( x2 & x5 ) | ( x2 & n18 ) | ( x5 & n18 ) ;
  assign n107 = ( x0 & x3 ) | ( x0 & n106 ) | ( x3 & n106 ) ;
  assign n108 = n18 & ~n107 ;
  assign n109 = ( n106 & ~n107 ) | ( n106 & n108 ) | ( ~n107 & n108 ) ;
  assign n110 = x4 & ~n109 ;
  assign n111 = x2 | x5 ;
  assign n112 = x3 | x5 ;
  assign n113 = x2 & ~n112 ;
  assign n114 = ( ~x2 & n111 ) | ( ~x2 & n113 ) | ( n111 & n113 ) ;
  assign n115 = x0 & n114 ;
  assign n116 = x4 | n115 ;
  assign n117 = ~n110 & n116 ;
  assign n118 = x1 & ~n117 ;
  assign n119 = ( x2 & x4 ) | ( x2 & x5 ) | ( x4 & x5 ) ;
  assign n120 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n121 = n119 & ~n120 ;
  assign n122 = x0 & n121 ;
  assign n123 = x1 | n122 ;
  assign n124 = ~n118 & n123 ;
  assign n125 = n105 | n124 ;
  assign n126 = ( n101 & ~n102 ) | ( n101 & n125 ) | ( ~n102 & n125 ) ;
  assign n127 = n96 | n126 ;
  assign n128 = ( n92 & ~n93 ) | ( n92 & n127 ) | ( ~n93 & n127 ) ;
  assign n129 = ( x2 & x3 ) | ( x2 & x4 ) | ( x3 & x4 ) ;
  assign n130 = x1 & ~n129 ;
  assign n131 = ~x1 & n129 ;
  assign n132 = n130 | n131 ;
  assign n133 = x5 & ~n132 ;
  assign n134 = ( ~x2 & n89 ) | ( ~x2 & n94 ) | ( n89 & n94 ) ;
  assign n135 = x4 & n134 ;
  assign n136 = x5 | n135 ;
  assign n137 = ~n133 & n136 ;
  assign n138 = ( x2 & x3 ) | ( x2 & x5 ) | ( x3 & x5 ) ;
  assign n139 = x3 & x4 ;
  assign n140 = ( x3 & x5 ) | ( x3 & n139 ) | ( x5 & n139 ) ;
  assign n141 = ( n37 & n138 ) | ( n37 & ~n140 ) | ( n138 & ~n140 ) ;
  assign n142 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n143 = ~x4 & n142 ;
  assign n144 = ( ~x3 & n142 ) | ( ~x3 & n143 ) | ( n142 & n143 ) ;
  assign y0 = n10 ;
  assign y1 = n16 ;
  assign y2 = n31 ;
  assign y3 = n59 ;
  assign y4 = n88 ;
  assign y5 = n128 ;
  assign y6 = n137 ;
  assign y7 = n141 ;
  assign y8 = n144 ;
  assign y9 = n71 ;
  assign y10 = 1'b0 ;
  assign y11 = x5 ;
endmodule
