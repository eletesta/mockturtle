module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 ;
  wire n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 ;
  assign n46 = ~x18 & x19 ;
  assign n47 = x21 & n46 ;
  assign n48 = x26 & n47 ;
  assign n49 = ~x29 & x30 ;
  assign n50 = ( x28 & n48 ) | ( x28 & n49 ) | ( n48 & n49 ) ;
  assign n51 = ~x28 & n50 ;
  assign n52 = ~x0 & x18 ;
  assign n53 = ~x20 & x21 ;
  assign n54 = ( x19 & n52 ) | ( x19 & n53 ) | ( n52 & n53 ) ;
  assign n55 = ~x19 & n54 ;
  assign n56 = ( x28 & n49 ) | ( x28 & n55 ) | ( n49 & n55 ) ;
  assign n57 = ~x28 & n56 ;
  assign n58 = x19 & x21 ;
  assign n59 = ( x20 & ~n52 ) | ( x20 & n58 ) | ( ~n52 & n58 ) ;
  assign n60 = n52 & n59 ;
  assign n61 = x24 & x30 ;
  assign n62 = ( x29 & n60 ) | ( x29 & n61 ) | ( n60 & n61 ) ;
  assign n63 = ~x29 & n62 ;
  assign n64 = x10 & x21 ;
  assign n65 = ( x18 & x19 ) | ( x18 & n64 ) | ( x19 & n64 ) ;
  assign n66 = ~x18 & n65 ;
  assign n67 = x25 & ~x29 ;
  assign n68 = ( x28 & n66 ) | ( x28 & n67 ) | ( n66 & n67 ) ;
  assign n69 = ~x28 & n68 ;
  assign n70 = x30 & n69 ;
  assign n71 = x24 & n47 ;
  assign n72 = ( x28 & n49 ) | ( x28 & n71 ) | ( n49 & n71 ) ;
  assign n73 = ~x28 & n72 ;
  assign n74 = ~x18 & x20 ;
  assign n75 = ( x0 & ~x19 ) | ( x0 & n74 ) | ( ~x19 & n74 ) ;
  assign n76 = ~x0 & n75 ;
  assign n77 = x21 & n76 ;
  assign n78 = ( x24 & x29 ) | ( x24 & n77 ) | ( x29 & n77 ) ;
  assign n79 = ~x29 & n78 ;
  assign n80 = x30 & n79 ;
  assign n81 = n73 | n80 ;
  assign n82 = n70 | n81 ;
  assign n83 = n63 | n82 ;
  assign n84 = ( ~n51 & n57 ) | ( ~n51 & n83 ) | ( n57 & n83 ) ;
  assign n85 = n51 | n84 ;
  assign n86 = n63 | n80 ;
  assign n87 = n51 | n70 ;
  assign n88 = n51 | n63 ;
  assign n89 = n73 | n88 ;
  assign n90 = ~x19 & x20 ;
  assign n91 = ( x0 & x18 ) | ( x0 & n90 ) | ( x18 & n90 ) ;
  assign n92 = ~x18 & n91 ;
  assign n93 = x21 & n92 ;
  assign n94 = ( x29 & n61 ) | ( x29 & n93 ) | ( n61 & n93 ) ;
  assign n95 = ~x29 & n94 ;
  assign n96 = x0 & x19 ;
  assign n97 = x18 & n96 ;
  assign n98 = x20 & n97 ;
  assign n99 = x21 & x30 ;
  assign n100 = ( x29 & n98 ) | ( x29 & n99 ) | ( n98 & n99 ) ;
  assign n101 = ~x29 & n100 ;
  assign n102 = x0 & ~x19 ;
  assign n103 = x18 & n102 ;
  assign n104 = ~x28 & n103 ;
  assign n105 = ( x20 & x21 ) | ( x20 & n104 ) | ( x21 & n104 ) ;
  assign n106 = ~x20 & n105 ;
  assign n107 = n49 & n106 ;
  assign n108 = x0 & x21 ;
  assign n109 = ( x18 & x19 ) | ( x18 & n108 ) | ( x19 & n108 ) ;
  assign n110 = ~x18 & n109 ;
  assign n111 = x28 & x30 ;
  assign n112 = ( x29 & n110 ) | ( x29 & n111 ) | ( n110 & n111 ) ;
  assign n113 = ~x29 & n112 ;
  assign n114 = n107 | n113 ;
  assign n115 = ( ~n95 & n101 ) | ( ~n95 & n114 ) | ( n101 & n114 ) ;
  assign n116 = n95 | n115 ;
  assign n117 = x10 & x18 ;
  assign n118 = ( x0 & x11 ) | ( x0 & n117 ) | ( x11 & n117 ) ;
  assign n119 = ~x11 & n118 ;
  assign n120 = x19 & ~x21 ;
  assign n121 = ( x20 & n119 ) | ( x20 & n120 ) | ( n119 & n120 ) ;
  assign n122 = ~x20 & n121 ;
  assign n123 = x25 & n122 ;
  assign n124 = ( x29 & x30 ) | ( x29 & n123 ) | ( x30 & n123 ) ;
  assign n125 = ~x30 & n124 ;
  assign n126 = x3 & x19 ;
  assign n127 = ( ~x0 & x18 ) | ( ~x0 & n126 ) | ( x18 & n126 ) ;
  assign n128 = x0 & n127 ;
  assign n129 = x20 & x27 ;
  assign n130 = ( x21 & n128 ) | ( x21 & n129 ) | ( n128 & n129 ) ;
  assign n131 = ~x21 & n130 ;
  assign n132 = ~x29 & n131 ;
  assign n133 = ~x30 & n132 ;
  assign n134 = x0 & ~x5 ;
  assign n135 = x19 & n134 ;
  assign n136 = x18 & n135 ;
  assign n137 = x20 & ~x27 ;
  assign n138 = ( x21 & n136 ) | ( x21 & n137 ) | ( n136 & n137 ) ;
  assign n139 = ~x21 & n138 ;
  assign n140 = x30 & n139 ;
  assign n141 = ( x28 & x29 ) | ( x28 & n140 ) | ( x29 & n140 ) ;
  assign n142 = ~x28 & n141 ;
  assign n143 = ~x4 & x19 ;
  assign n144 = ( x0 & x18 ) | ( x0 & n143 ) | ( x18 & n143 ) ;
  assign n145 = ~x0 & n144 ;
  assign n146 = ( x21 & n137 ) | ( x21 & n145 ) | ( n137 & n145 ) ;
  assign n147 = ~x21 & n146 ;
  assign n148 = x28 & n147 ;
  assign n149 = ( x29 & x30 ) | ( x29 & n148 ) | ( x30 & n148 ) ;
  assign n150 = ~x30 & n149 ;
  assign n151 = n142 | n150 ;
  assign n152 = n133 | n151 ;
  assign n153 = ~x21 & x26 ;
  assign n154 = ( x20 & n97 ) | ( x20 & n153 ) | ( n97 & n153 ) ;
  assign n155 = ~x20 & n154 ;
  assign n156 = ~x30 & n155 ;
  assign n157 = ( x28 & x29 ) | ( x28 & n156 ) | ( x29 & n156 ) ;
  assign n158 = ~x28 & n157 ;
  assign n159 = x11 & x19 ;
  assign n160 = ( ~x0 & x18 ) | ( ~x0 & n159 ) | ( x18 & n159 ) ;
  assign n161 = x0 & n160 ;
  assign n162 = ( x20 & n153 ) | ( x20 & n161 ) | ( n153 & n161 ) ;
  assign n163 = ~x20 & n162 ;
  assign n164 = ( x29 & n111 ) | ( x29 & n163 ) | ( n111 & n163 ) ;
  assign n165 = ~x29 & n164 ;
  assign n166 = ( x11 & x18 ) | ( x11 & n96 ) | ( x18 & n96 ) ;
  assign n167 = ~x11 & n166 ;
  assign n168 = ( x20 & n153 ) | ( x20 & n167 ) | ( n153 & n167 ) ;
  assign n169 = ~x20 & n168 ;
  assign n170 = ( x29 & n111 ) | ( x29 & n169 ) | ( n111 & n169 ) ;
  assign n171 = ~x29 & n170 ;
  assign n172 = n165 | n171 ;
  assign n173 = n158 | n172 ;
  assign n174 = ( ~n125 & n152 ) | ( ~n125 & n173 ) | ( n152 & n173 ) ;
  assign n175 = n125 | n174 ;
  assign n176 = x0 & ~x3 ;
  assign n177 = ( x2 & ~x18 ) | ( x2 & n176 ) | ( ~x18 & n176 ) ;
  assign n178 = ~x2 & n177 ;
  assign n179 = ~x21 & n178 ;
  assign n180 = ( x19 & x20 ) | ( x19 & n179 ) | ( x20 & n179 ) ;
  assign n181 = ~x19 & n180 ;
  assign n182 = ( x29 & n111 ) | ( x29 & n181 ) | ( n111 & n181 ) ;
  assign n183 = ~x29 & n182 ;
  assign n184 = ~x28 & n92 ;
  assign n185 = ( x21 & x23 ) | ( x21 & n184 ) | ( x23 & n184 ) ;
  assign n186 = ~x21 & n185 ;
  assign n187 = ~x30 & n186 ;
  assign n188 = x29 & n187 ;
  assign n189 = x2 & ~x18 ;
  assign n190 = ( x0 & x3 ) | ( x0 & n189 ) | ( x3 & n189 ) ;
  assign n191 = ~x3 & n190 ;
  assign n192 = ~x20 & n191 ;
  assign n193 = ( x19 & ~x21 ) | ( x19 & n192 ) | ( ~x21 & n192 ) ;
  assign n194 = ~x19 & n193 ;
  assign n195 = ( x29 & n111 ) | ( x29 & n194 ) | ( n111 & n194 ) ;
  assign n196 = ~x29 & n195 ;
  assign n197 = ~x15 & n134 ;
  assign n198 = x11 & n197 ;
  assign n199 = x18 & x20 ;
  assign n200 = ( x19 & n198 ) | ( x19 & n199 ) | ( n198 & n199 ) ;
  assign n201 = ~x19 & n200 ;
  assign n202 = x21 & n201 ;
  assign n203 = ( x26 & x28 ) | ( x26 & n202 ) | ( x28 & n202 ) ;
  assign n204 = ~x28 & n203 ;
  assign n205 = n49 & n204 ;
  assign n206 = ~x11 & n134 ;
  assign n207 = ~x15 & n206 ;
  assign n208 = ( x19 & n199 ) | ( x19 & n207 ) | ( n199 & n207 ) ;
  assign n209 = ~x19 & n208 ;
  assign n210 = x21 & n209 ;
  assign n211 = ( x26 & x28 ) | ( x26 & n210 ) | ( x28 & n210 ) ;
  assign n212 = ~x28 & n211 ;
  assign n213 = n49 & n212 ;
  assign n214 = x11 & n134 ;
  assign n215 = x10 & n214 ;
  assign n216 = ~x19 & n215 ;
  assign n217 = ( x15 & x18 ) | ( x15 & n216 ) | ( x18 & n216 ) ;
  assign n218 = ~x15 & n217 ;
  assign n219 = x20 & x25 ;
  assign n220 = ( x21 & ~n218 ) | ( x21 & n219 ) | ( ~n218 & n219 ) ;
  assign n221 = n218 & n220 ;
  assign n222 = ( x28 & n49 ) | ( x28 & n221 ) | ( n49 & n221 ) ;
  assign n223 = ~x28 & n222 ;
  assign n224 = ( x3 & ~x18 ) | ( x3 & n134 ) | ( ~x18 & n134 ) ;
  assign n225 = ~x3 & n224 ;
  assign n226 = ~x20 & n225 ;
  assign n227 = ( x19 & ~x21 ) | ( x19 & n226 ) | ( ~x21 & n226 ) ;
  assign n228 = ~x19 & n227 ;
  assign n229 = ~x30 & n228 ;
  assign n230 = ( x28 & x29 ) | ( x28 & n229 ) | ( x29 & n229 ) ;
  assign n231 = ~x28 & n230 ;
  assign n232 = n223 | n231 ;
  assign n233 = ( ~n205 & n213 ) | ( ~n205 & n232 ) | ( n213 & n232 ) ;
  assign n234 = n205 | n233 ;
  assign n235 = n196 | n234 ;
  assign n236 = ( ~n183 & n188 ) | ( ~n183 & n235 ) | ( n188 & n235 ) ;
  assign n237 = n183 | n236 ;
  assign n238 = x22 & x30 ;
  assign n239 = ( x29 & n93 ) | ( x29 & n238 ) | ( n93 & n238 ) ;
  assign n240 = ~x29 & n239 ;
  assign n241 = x10 & ~x18 ;
  assign n242 = ( x0 & x11 ) | ( x0 & n241 ) | ( x11 & n241 ) ;
  assign n243 = ~x11 & n242 ;
  assign n244 = x21 & n243 ;
  assign n245 = ( x19 & x20 ) | ( x19 & n244 ) | ( x20 & n244 ) ;
  assign n246 = ~x19 & n245 ;
  assign n247 = x25 & x30 ;
  assign n248 = ( x29 & n246 ) | ( x29 & n247 ) | ( n246 & n247 ) ;
  assign n249 = ~x29 & n248 ;
  assign n250 = n240 | n249 ;
  assign n251 = x11 & ~x19 ;
  assign n252 = ( x0 & x18 ) | ( x0 & n251 ) | ( x18 & n251 ) ;
  assign n253 = ~x18 & n252 ;
  assign n254 = x20 & x26 ;
  assign n255 = ( x21 & ~n253 ) | ( x21 & n254 ) | ( ~n253 & n254 ) ;
  assign n256 = n253 & n255 ;
  assign n257 = n49 & n256 ;
  assign n258 = ( x15 & n46 ) | ( x15 & n134 ) | ( n46 & n134 ) ;
  assign n259 = ~x15 & n258 ;
  assign n260 = x20 & x22 ;
  assign n261 = ( x21 & ~n259 ) | ( x21 & n260 ) | ( ~n259 & n260 ) ;
  assign n262 = n259 & n261 ;
  assign n263 = ( x28 & n49 ) | ( x28 & n262 ) | ( n49 & n262 ) ;
  assign n264 = ~x28 & n263 ;
  assign n265 = x10 & n206 ;
  assign n266 = ~x19 & n265 ;
  assign n267 = ( x15 & x18 ) | ( x15 & n266 ) | ( x18 & n266 ) ;
  assign n268 = ~x15 & n267 ;
  assign n269 = ( x21 & n219 ) | ( x21 & ~n268 ) | ( n219 & ~n268 ) ;
  assign n270 = n268 & n269 ;
  assign n271 = ( x28 & n49 ) | ( x28 & n270 ) | ( n49 & n270 ) ;
  assign n272 = ~x28 & n271 ;
  assign n273 = ~x19 & n134 ;
  assign n274 = ( x15 & x18 ) | ( x15 & n273 ) | ( x18 & n273 ) ;
  assign n275 = ~x15 & n274 ;
  assign n276 = ( x21 & n260 ) | ( x21 & ~n275 ) | ( n260 & ~n275 ) ;
  assign n277 = n275 & n276 ;
  assign n278 = ( x28 & n49 ) | ( x28 & n277 ) | ( n49 & n277 ) ;
  assign n279 = ~x28 & n278 ;
  assign n280 = n272 | n279 ;
  assign n281 = n264 | n280 ;
  assign n282 = n257 | n281 ;
  assign n283 = x0 & x10 ;
  assign n284 = ( x11 & x18 ) | ( x11 & n283 ) | ( x18 & n283 ) ;
  assign n285 = ~x18 & n284 ;
  assign n286 = x21 & n285 ;
  assign n287 = ( x19 & x20 ) | ( x19 & n286 ) | ( x20 & n286 ) ;
  assign n288 = ~x19 & n287 ;
  assign n289 = ( x29 & n247 ) | ( x29 & n288 ) | ( n247 & n288 ) ;
  assign n290 = ~x29 & n289 ;
  assign n291 = x0 & ~x18 ;
  assign n292 = ( x11 & ~x19 ) | ( x11 & n291 ) | ( ~x19 & n291 ) ;
  assign n293 = ~x11 & n292 ;
  assign n294 = ( x21 & n254 ) | ( x21 & ~n293 ) | ( n254 & ~n293 ) ;
  assign n295 = n293 & n294 ;
  assign n296 = n49 & n295 ;
  assign n297 = n290 | n296 ;
  assign n298 = n282 | n297 ;
  assign n299 = ( ~n237 & n250 ) | ( ~n237 & n298 ) | ( n250 & n298 ) ;
  assign n300 = n237 | n299 ;
  assign n301 = ~x21 & x22 ;
  assign n302 = ( x20 & n97 ) | ( x20 & n301 ) | ( n97 & n301 ) ;
  assign n303 = ~x20 & n302 ;
  assign n304 = ~x30 & n303 ;
  assign n305 = x29 & n304 ;
  assign n306 = x0 & x20 ;
  assign n307 = ( x18 & x19 ) | ( x18 & n306 ) | ( x19 & n306 ) ;
  assign n308 = ~x18 & n307 ;
  assign n309 = n301 & n308 ;
  assign n310 = x28 & n309 ;
  assign n311 = ( x29 & x30 ) | ( x29 & n310 ) | ( x30 & n310 ) ;
  assign n312 = ~x30 & n311 ;
  assign n313 = n46 & n134 ;
  assign n314 = ( x21 & n260 ) | ( x21 & n313 ) | ( n260 & n313 ) ;
  assign n315 = ~x21 & n314 ;
  assign n316 = ~x30 & n315 ;
  assign n317 = ( x28 & x29 ) | ( x28 & n316 ) | ( x29 & n316 ) ;
  assign n318 = ~x28 & n317 ;
  assign n319 = x0 & x17 ;
  assign n320 = ( x18 & x19 ) | ( x18 & n319 ) | ( x19 & n319 ) ;
  assign n321 = ~x19 & n320 ;
  assign n322 = ( x21 & n254 ) | ( x21 & n321 ) | ( n254 & n321 ) ;
  assign n323 = ~x21 & n322 ;
  assign n324 = ~x30 & n323 ;
  assign n325 = ( x28 & x29 ) | ( x28 & n324 ) | ( x29 & n324 ) ;
  assign n326 = ~x28 & n325 ;
  assign n327 = ( x17 & x18 ) | ( x17 & n102 ) | ( x18 & n102 ) ;
  assign n328 = ~x17 & n327 ;
  assign n329 = ( x21 & n254 ) | ( x21 & n328 ) | ( n254 & n328 ) ;
  assign n330 = ~x21 & n329 ;
  assign n331 = ~x30 & n330 ;
  assign n332 = ( x28 & x29 ) | ( x28 & n331 ) | ( x29 & n331 ) ;
  assign n333 = ~x28 & n332 ;
  assign n334 = n326 | n333 ;
  assign n335 = n318 | n334 ;
  assign n336 = n312 | n335 ;
  assign n337 = ( ~x0 & x11 ) | ( ~x0 & n117 ) | ( x11 & n117 ) ;
  assign n338 = x0 & n337 ;
  assign n339 = ( x20 & n120 ) | ( x20 & n338 ) | ( n120 & n338 ) ;
  assign n340 = ~x20 & n339 ;
  assign n341 = x25 & n340 ;
  assign n342 = ( x29 & x30 ) | ( x29 & n341 ) | ( x30 & n341 ) ;
  assign n343 = ~x30 & n342 ;
  assign n344 = ( x11 & x18 ) | ( x11 & n102 ) | ( x18 & n102 ) ;
  assign n345 = ~x11 & n344 ;
  assign n346 = ( x21 & n254 ) | ( x21 & n345 ) | ( n254 & n345 ) ;
  assign n347 = ~x21 & n346 ;
  assign n348 = ( x29 & n111 ) | ( x29 & n347 ) | ( n111 & n347 ) ;
  assign n349 = ~x29 & n348 ;
  assign n350 = x0 & x11 ;
  assign n351 = ( x18 & x19 ) | ( x18 & n350 ) | ( x19 & n350 ) ;
  assign n352 = ~x19 & n351 ;
  assign n353 = ( x21 & n254 ) | ( x21 & n352 ) | ( n254 & n352 ) ;
  assign n354 = ~x21 & n353 ;
  assign n355 = ( x29 & n111 ) | ( x29 & n354 ) | ( n111 & n354 ) ;
  assign n356 = ~x29 & n355 ;
  assign n357 = n349 | n356 ;
  assign n358 = n343 | n357 ;
  assign n359 = ( ~n305 & n336 ) | ( ~n305 & n358 ) | ( n336 & n358 ) ;
  assign n360 = n305 | n359 ;
  assign n361 = n300 | n360 ;
  assign n362 = n175 | n361 ;
  assign n363 = n272 | n290 ;
  assign n364 = n249 | n363 ;
  assign n365 = n125 | n364 ;
  assign n366 = ( ~n223 & n343 ) | ( ~n223 & n365 ) | ( n343 & n365 ) ;
  assign n367 = n223 | n366 ;
  assign n368 = n250 | n264 ;
  assign n369 = n296 | n368 ;
  assign n370 = n231 | n280 ;
  assign n371 = ( ~n213 & n369 ) | ( ~n213 & n370 ) | ( n369 & n370 ) ;
  assign n372 = n213 | n371 ;
  assign n373 = n183 | n356 ;
  assign n374 = ( ~n305 & n312 ) | ( ~n305 & n373 ) | ( n312 & n373 ) ;
  assign n375 = n305 | n374 ;
  assign n376 = n171 | n375 ;
  assign n377 = ( n125 & ~n150 ) | ( n125 & n376 ) | ( ~n150 & n376 ) ;
  assign n378 = n150 | n377 ;
  assign n379 = n372 | n378 ;
  assign n380 = n133 | n188 ;
  assign n381 = n196 | n380 ;
  assign n382 = ~x19 & x21 ;
  assign n383 = ( x18 & ~x20 ) | ( x18 & n382 ) | ( ~x20 & n382 ) ;
  assign n384 = ~x18 & n383 ;
  assign n385 = x22 & x29 ;
  assign n386 = ( x28 & n384 ) | ( x28 & n385 ) | ( n384 & n385 ) ;
  assign n387 = ~x28 & n386 ;
  assign n388 = x30 & n387 ;
  assign n389 = x18 | x20 ;
  assign n390 = ( ~x9 & x19 ) | ( ~x9 & n389 ) | ( x19 & n389 ) ;
  assign n391 = x9 | n390 ;
  assign n392 = x21 & ~n391 ;
  assign n393 = ( x22 & x28 ) | ( x22 & n392 ) | ( x28 & n392 ) ;
  assign n394 = ~x28 & n393 ;
  assign n395 = ~x30 & n394 ;
  assign n396 = x29 & n395 ;
  assign n397 = ~x38 & n396 ;
  assign n398 = ~x39 & n397 ;
  assign n399 = ~x41 & n398 ;
  assign n400 = ( x40 & ~x42 ) | ( x40 & n399 ) | ( ~x42 & n399 ) ;
  assign n401 = ~x40 & n400 ;
  assign n402 = ~x43 & x44 ;
  assign n403 = n401 & n402 ;
  assign n404 = x39 & x42 ;
  assign n405 = ( x41 & n397 ) | ( x41 & n404 ) | ( n397 & n404 ) ;
  assign n406 = ~x41 & n405 ;
  assign n407 = ~x41 & x42 ;
  assign n408 = n398 & n407 ;
  assign n409 = x39 & ~x42 ;
  assign n410 = ( x41 & n397 ) | ( x41 & n409 ) | ( n397 & n409 ) ;
  assign n411 = ~x41 & n410 ;
  assign n412 = n408 | n411 ;
  assign n413 = n406 | n412 ;
  assign n414 = n403 | n413 ;
  assign n415 = n388 | n414 ;
  assign n416 = ( x17 & x19 ) | ( x17 & n199 ) | ( x19 & n199 ) ;
  assign n417 = ~x19 & n416 ;
  assign n418 = n153 & n417 ;
  assign n419 = ~x28 & n418 ;
  assign n420 = ~x30 & n419 ;
  assign n421 = x29 & n420 ;
  assign n422 = ( x17 & x18 ) | ( x17 & n90 ) | ( x18 & n90 ) ;
  assign n423 = ~x17 & n422 ;
  assign n424 = ~x28 & n423 ;
  assign n425 = ( x21 & x26 ) | ( x21 & n424 ) | ( x26 & n424 ) ;
  assign n426 = ~x21 & n425 ;
  assign n427 = x30 & n426 ;
  assign n428 = x29 & n427 ;
  assign n429 = x18 & ~x21 ;
  assign n430 = ( x19 & x20 ) | ( x19 & n429 ) | ( x20 & n429 ) ;
  assign n431 = ~x19 & n430 ;
  assign n432 = x26 & x29 ;
  assign n433 = ( x28 & ~n431 ) | ( x28 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = n431 & n433 ;
  assign n435 = ~x30 & n434 ;
  assign n436 = ~x21 & n46 ;
  assign n437 = x20 & n436 ;
  assign n438 = ~x28 & n437 ;
  assign n439 = x22 & n438 ;
  assign n440 = x30 & n439 ;
  assign n441 = x29 & n440 ;
  assign n442 = x28 & n437 ;
  assign n443 = x22 & n442 ;
  assign n444 = x30 & n443 ;
  assign n445 = x29 & n444 ;
  assign n446 = x1 & ~x20 ;
  assign n447 = ( x18 & x19 ) | ( x18 & n446 ) | ( x19 & n446 ) ;
  assign n448 = ~x18 & n447 ;
  assign n449 = ~x21 & n448 ;
  assign n450 = x23 & n449 ;
  assign n451 = ( x29 & x30 ) | ( x29 & n450 ) | ( x30 & n450 ) ;
  assign n452 = ~x30 & n451 ;
  assign n453 = n445 | n452 ;
  assign n454 = n441 | n453 ;
  assign n455 = n435 | n454 ;
  assign n456 = ( ~n421 & n428 ) | ( ~n421 & n455 ) | ( n428 & n455 ) ;
  assign n457 = n421 | n456 ;
  assign n458 = x41 & n397 ;
  assign n459 = x38 & n396 ;
  assign n460 = x9 & ~x19 ;
  assign n461 = ( x18 & ~x20 ) | ( x18 & n460 ) | ( ~x20 & n460 ) ;
  assign n462 = ~x18 & n461 ;
  assign n463 = x21 & n462 ;
  assign n464 = ( x22 & x28 ) | ( x22 & n463 ) | ( x28 & n463 ) ;
  assign n465 = ~x28 & n464 ;
  assign n466 = n49 & n465 ;
  assign n467 = ~x33 & x39 ;
  assign n468 = ( x31 & n466 ) | ( x31 & n467 ) | ( n466 & n467 ) ;
  assign n469 = ~x31 & n468 ;
  assign n470 = x18 & x19 ;
  assign n471 = ( x20 & x21 ) | ( x20 & n470 ) | ( x21 & n470 ) ;
  assign n472 = ~x21 & n471 ;
  assign n473 = x29 & n472 ;
  assign n474 = ( x27 & x28 ) | ( x27 & n473 ) | ( x28 & n473 ) ;
  assign n475 = ~x27 & n474 ;
  assign n476 = x30 & n475 ;
  assign n477 = n49 & n394 ;
  assign n478 = x27 & x30 ;
  assign n479 = ( x29 & n472 ) | ( x29 & n478 ) | ( n472 & n478 ) ;
  assign n480 = ~x29 & n479 ;
  assign n481 = n477 | n480 ;
  assign n482 = n476 | n481 ;
  assign n483 = n469 | n482 ;
  assign n484 = ( ~n458 & n459 ) | ( ~n458 & n483 ) | ( n459 & n483 ) ;
  assign n485 = n458 | n484 ;
  assign n486 = ~x29 & n472 ;
  assign n487 = ( x27 & x28 ) | ( x27 & n486 ) | ( x28 & n486 ) ;
  assign n488 = ~x27 & n487 ;
  assign n489 = ~x30 & n488 ;
  assign n490 = ( x18 & x20 ) | ( x18 & n120 ) | ( x20 & n120 ) ;
  assign n491 = ~x20 & n490 ;
  assign n492 = x28 & n491 ;
  assign n493 = x26 & n492 ;
  assign n494 = ~x30 & n493 ;
  assign n495 = x29 & n494 ;
  assign n496 = ( x29 & n238 ) | ( x29 & ~n491 ) | ( n238 & ~n491 ) ;
  assign n497 = n491 & n496 ;
  assign n498 = ~x28 & n491 ;
  assign n499 = x26 & n498 ;
  assign n500 = x30 & n499 ;
  assign n501 = x29 & n500 ;
  assign n502 = ( x29 & n247 ) | ( x29 & ~n491 ) | ( n247 & ~n491 ) ;
  assign n503 = n491 & n502 ;
  assign n504 = n501 | n503 ;
  assign n505 = n497 | n504 ;
  assign n506 = n495 | n505 ;
  assign n507 = n489 | n506 ;
  assign n508 = n485 | n507 ;
  assign n509 = ( ~n415 & n457 ) | ( ~n415 & n508 ) | ( n457 & n508 ) ;
  assign n510 = n415 | n509 ;
  assign n511 = ( ~x18 & x20 ) | ( ~x18 & n58 ) | ( x20 & n58 ) ;
  assign n512 = x18 & n511 ;
  assign n513 = ~x30 & n512 ;
  assign n514 = x29 & n513 ;
  assign n515 = x25 & x29 ;
  assign n516 = ( x11 & x19 ) | ( x11 & n199 ) | ( x19 & n199 ) ;
  assign n517 = ~x19 & n516 ;
  assign n518 = x21 & n517 ;
  assign n519 = ( x28 & n515 ) | ( x28 & n518 ) | ( n515 & n518 ) ;
  assign n520 = ~x28 & n519 ;
  assign n521 = ( x11 & x18 ) | ( x11 & n90 ) | ( x18 & n90 ) ;
  assign n522 = ~x11 & n521 ;
  assign n523 = x21 & n522 ;
  assign n524 = ( x28 & n432 ) | ( x28 & n523 ) | ( n432 & n523 ) ;
  assign n525 = ~x28 & n524 ;
  assign n526 = x30 & ~n525 ;
  assign n527 = ( n520 & n525 ) | ( n520 & ~n526 ) | ( n525 & ~n526 ) ;
  assign n528 = ( x28 & n432 ) | ( x28 & n518 ) | ( n432 & n518 ) ;
  assign n529 = ~x28 & n528 ;
  assign n530 = x22 & n449 ;
  assign n531 = ( x29 & x30 ) | ( x29 & n530 ) | ( x30 & n530 ) ;
  assign n532 = ~x30 & n531 ;
  assign n533 = ( x18 & ~x21 ) | ( x18 & n90 ) | ( ~x21 & n90 ) ;
  assign n534 = ~x18 & n533 ;
  assign n535 = x30 & n534 ;
  assign n536 = ( x28 & x29 ) | ( x28 & n535 ) | ( x29 & n535 ) ;
  assign n537 = ~x28 & n536 ;
  assign n538 = x28 & n534 ;
  assign n539 = ( x29 & x30 ) | ( x29 & n538 ) | ( x30 & n538 ) ;
  assign n540 = ~x30 & n539 ;
  assign n541 = x19 | x21 ;
  assign n542 = ( ~x18 & x20 ) | ( ~x18 & n541 ) | ( x20 & n541 ) ;
  assign n543 = x18 | n542 ;
  assign n544 = x30 & ~n543 ;
  assign n545 = ( x28 & x29 ) | ( x28 & n544 ) | ( x29 & n544 ) ;
  assign n546 = ~x28 & n545 ;
  assign n547 = x28 & ~n543 ;
  assign n548 = ( x29 & x30 ) | ( x29 & n547 ) | ( x30 & n547 ) ;
  assign n549 = ~x30 & n548 ;
  assign n550 = n546 | n549 ;
  assign n551 = n540 | n550 ;
  assign n552 = ( ~n532 & n537 ) | ( ~n532 & n551 ) | ( n537 & n551 ) ;
  assign n553 = n532 | n552 ;
  assign n554 = n529 | n553 ;
  assign n555 = ( ~n514 & n527 ) | ( ~n514 & n554 ) | ( n527 & n554 ) ;
  assign n556 = n514 | n555 ;
  assign n557 = x20 & n47 ;
  assign n558 = ( x28 & n385 ) | ( x28 & n557 ) | ( n385 & n557 ) ;
  assign n559 = ~x28 & n558 ;
  assign n560 = ~x30 & n559 ;
  assign n561 = ( x18 & x19 ) | ( x18 & n53 ) | ( x19 & n53 ) ;
  assign n562 = ~x19 & n561 ;
  assign n563 = ~x30 & n562 ;
  assign n564 = ( x28 & x29 ) | ( x28 & n563 ) | ( x29 & n563 ) ;
  assign n565 = ~x28 & n564 ;
  assign n566 = x28 & n47 ;
  assign n567 = ( x29 & x30 ) | ( x29 & n566 ) | ( x30 & n566 ) ;
  assign n568 = ~x30 & n567 ;
  assign n569 = ( x28 & n515 ) | ( x28 & n523 ) | ( n515 & n523 ) ;
  assign n570 = ~x28 & n569 ;
  assign n571 = ~x30 & n570 ;
  assign n572 = x18 & x21 ;
  assign n573 = ( x19 & x20 ) | ( x19 & n572 ) | ( x20 & n572 ) ;
  assign n574 = ~x19 & n573 ;
  assign n575 = ( x28 & n385 ) | ( x28 & n574 ) | ( n385 & n574 ) ;
  assign n576 = ~x28 & n575 ;
  assign n577 = ~x30 & n576 ;
  assign n578 = n571 | n577 ;
  assign n579 = n568 | n578 ;
  assign n580 = ( ~n560 & n565 ) | ( ~n560 & n579 ) | ( n565 & n579 ) ;
  assign n581 = n560 | n580 ;
  assign n582 = x21 & n448 ;
  assign n583 = ( x23 & x28 ) | ( x23 & n582 ) | ( x28 & n582 ) ;
  assign n584 = ~x28 & n583 ;
  assign n585 = n49 & n584 ;
  assign n586 = ( x18 & x20 ) | ( x18 & n382 ) | ( x20 & n382 ) ;
  assign n587 = ~x18 & n586 ;
  assign n588 = ~x30 & n587 ;
  assign n589 = ( x26 & x29 ) | ( x26 & n588 ) | ( x29 & n588 ) ;
  assign n590 = ~x26 & n589 ;
  assign n591 = x26 & n587 ;
  assign n592 = ( x29 & x30 ) | ( x29 & n591 ) | ( x30 & n591 ) ;
  assign n593 = ~x30 & n592 ;
  assign n594 = n590 | n593 ;
  assign n595 = x26 & x30 ;
  assign n596 = ( x29 & ~n587 ) | ( x29 & n595 ) | ( ~n587 & n595 ) ;
  assign n597 = n587 & n596 ;
  assign n598 = ( x22 & x28 ) | ( x22 & n582 ) | ( x28 & n582 ) ;
  assign n599 = ~x28 & n598 ;
  assign n600 = n49 & n599 ;
  assign n601 = x24 & n587 ;
  assign n602 = ( x29 & x30 ) | ( x29 & n601 ) | ( x30 & n601 ) ;
  assign n603 = ~x30 & n602 ;
  assign n604 = n600 | n603 ;
  assign n605 = n597 | n604 ;
  assign n606 = ( ~n585 & n594 ) | ( ~n585 & n605 ) | ( n594 & n605 ) ;
  assign n607 = n585 | n606 ;
  assign n608 = n581 | n607 ;
  assign n609 = ( ~n510 & n556 ) | ( ~n510 & n608 ) | ( n556 & n608 ) ;
  assign n610 = n510 | n609 ;
  assign n611 = ~x44 & n401 ;
  assign n612 = x43 & n611 ;
  assign n613 = ( x3 & x19 ) | ( x3 & n199 ) | ( x19 & n199 ) ;
  assign n614 = ~x3 & n613 ;
  assign n615 = ~x29 & n614 ;
  assign n616 = ( x21 & x27 ) | ( x21 & n615 ) | ( x27 & n615 ) ;
  assign n617 = ~x21 & n616 ;
  assign n618 = ~x30 & n617 ;
  assign n619 = n489 | n618 ;
  assign n620 = x28 & ~x30 ;
  assign n621 = ( x29 & n418 ) | ( x29 & n620 ) | ( n418 & n620 ) ;
  assign n622 = ~x29 & n621 ;
  assign n623 = ~x29 & n493 ;
  assign n624 = ~x30 & n623 ;
  assign n625 = n501 | n624 ;
  assign n626 = n441 | n625 ;
  assign n627 = ( ~n421 & n622 ) | ( ~n421 & n626 ) | ( n622 & n626 ) ;
  assign n628 = n421 | n627 ;
  assign n629 = n480 | n628 ;
  assign n630 = ( ~n612 & n619 ) | ( ~n612 & n629 ) | ( n619 & n629 ) ;
  assign n631 = n612 | n630 ;
  assign n632 = n514 | n546 ;
  assign n633 = n549 | n632 ;
  assign n634 = n540 | n633 ;
  assign n635 = n537 | n634 ;
  assign n636 = x30 & n559 ;
  assign n637 = ( x29 & ~n47 ) | ( x29 & n111 ) | ( ~n47 & n111 ) ;
  assign n638 = n47 & n637 ;
  assign n639 = n560 | n638 ;
  assign n640 = n568 | n639 ;
  assign n641 = x30 & n562 ;
  assign n642 = ( x28 & x29 ) | ( x28 & n641 ) | ( x29 & n641 ) ;
  assign n643 = ~x28 & n642 ;
  assign n644 = n570 | n576 ;
  assign n645 = n643 | n644 ;
  assign n646 = n565 | n645 ;
  assign n647 = ( ~n636 & n640 ) | ( ~n636 & n646 ) | ( n640 & n646 ) ;
  assign n648 = n636 | n647 ;
  assign n649 = n597 | n603 ;
  assign n650 = x23 & n46 ;
  assign n651 = ( x20 & x21 ) | ( x20 & n650 ) | ( x21 & n650 ) ;
  assign n652 = ~x20 & n651 ;
  assign n653 = ~x30 & n652 ;
  assign n654 = ( x28 & x29 ) | ( x28 & n653 ) | ( x29 & n653 ) ;
  assign n655 = ~x28 & n654 ;
  assign n656 = x22 & n46 ;
  assign n657 = ( x20 & x21 ) | ( x20 & n656 ) | ( x21 & n656 ) ;
  assign n658 = ~x20 & n657 ;
  assign n659 = ~x30 & n658 ;
  assign n660 = ( x28 & x29 ) | ( x28 & n659 ) | ( x29 & n659 ) ;
  assign n661 = ~x28 & n660 ;
  assign n662 = ( x29 & n61 ) | ( x29 & ~n587 ) | ( n61 & ~n587 ) ;
  assign n663 = n587 & n662 ;
  assign n664 = n600 | n663 ;
  assign n665 = n661 | n664 ;
  assign n666 = ( ~n585 & n655 ) | ( ~n585 & n665 ) | ( n655 & n665 ) ;
  assign n667 = n585 | n666 ;
  assign n668 = x30 & n587 ;
  assign n669 = ( x26 & x29 ) | ( x26 & n668 ) | ( x29 & n668 ) ;
  assign n670 = ~x26 & n669 ;
  assign n671 = n590 | n670 ;
  assign n672 = n593 | n671 ;
  assign n673 = n667 | n672 ;
  assign n674 = ( ~n648 & n649 ) | ( ~n648 & n673 ) | ( n649 & n673 ) ;
  assign n675 = n648 | n674 ;
  assign n676 = ~x30 & n520 ;
  assign n677 = n525 | n529 ;
  assign n678 = ( n520 & ~n676 ) | ( n520 & n677 ) | ( ~n676 & n677 ) ;
  assign n679 = n675 | n678 ;
  assign n680 = ( ~n631 & n635 ) | ( ~n631 & n679 ) | ( n635 & n679 ) ;
  assign n681 = n631 | n680 ;
  assign n682 = n476 | n618 ;
  assign n683 = n435 | n503 ;
  assign n684 = ( n497 & ~n501 ) | ( n497 & n683 ) | ( ~n501 & n683 ) ;
  assign n685 = n501 | n684 ;
  assign n686 = n495 | n624 ;
  assign n687 = n489 | n686 ;
  assign n688 = n685 | n687 ;
  assign n689 = ~x43 & n401 ;
  assign n690 = ~x44 & n689 ;
  assign n691 = n403 | n477 ;
  assign n692 = n690 | n691 ;
  assign n693 = n688 | n692 ;
  assign n694 = ( ~n480 & n682 ) | ( ~n480 & n693 ) | ( n682 & n693 ) ;
  assign n695 = n480 | n694 ;
  assign n696 = n428 | n454 ;
  assign n697 = ( ~n421 & n622 ) | ( ~n421 & n696 ) | ( n622 & n696 ) ;
  assign n698 = n421 | n697 ;
  assign n699 = x30 & n520 ;
  assign n700 = x30 & n570 ;
  assign n701 = n676 | n700 ;
  assign n702 = x30 & n576 ;
  assign n703 = n571 | n702 ;
  assign n704 = n577 | n643 ;
  assign n705 = n703 | n704 ;
  assign n706 = ( ~n699 & n701 ) | ( ~n699 & n705 ) | ( n701 & n705 ) ;
  assign n707 = n699 | n706 ;
  assign n708 = n568 | n655 ;
  assign n709 = n638 | n708 ;
  assign n710 = n636 | n709 ;
  assign n711 = ( ~n560 & n565 ) | ( ~n560 & n710 ) | ( n565 & n710 ) ;
  assign n712 = n560 | n711 ;
  assign n713 = x30 & n529 ;
  assign n714 = ( x19 & x20 ) | ( x19 & n117 ) | ( x20 & n117 ) ;
  assign n715 = ~x20 & n714 ;
  assign n716 = ( x25 & n99 ) | ( x25 & ~n715 ) | ( n99 & ~n715 ) ;
  assign n717 = n715 & n716 ;
  assign n718 = ( x18 & x20 ) | ( x18 & n58 ) | ( x20 & n58 ) ;
  assign n719 = ~x20 & n718 ;
  assign n720 = x30 & n719 ;
  assign n721 = x26 & n720 ;
  assign n722 = ( n525 & ~n526 ) | ( n525 & n529 ) | ( ~n526 & n529 ) ;
  assign n723 = n721 | n722 ;
  assign n724 = ( ~n713 & n717 ) | ( ~n713 & n723 ) | ( n717 & n723 ) ;
  assign n725 = n713 | n724 ;
  assign n726 = x29 & n587 ;
  assign n727 = n603 | n726 ;
  assign n728 = ( ~n661 & n663 ) | ( ~n661 & n727 ) | ( n663 & n727 ) ;
  assign n729 = n661 | n728 ;
  assign n730 = n725 | n729 ;
  assign n731 = ( ~n707 & n712 ) | ( ~n707 & n730 ) | ( n712 & n730 ) ;
  assign n732 = n707 | n731 ;
  assign n733 = x30 & n512 ;
  assign n734 = x29 & n733 ;
  assign n735 = n514 | n550 ;
  assign n736 = n734 | n735 ;
  assign n737 = n540 | n736 ;
  assign n738 = ( ~n532 & n537 ) | ( ~n532 & n737 ) | ( n537 & n737 ) ;
  assign n739 = n532 | n738 ;
  assign n740 = n732 | n739 ;
  assign n741 = ( ~n695 & n698 ) | ( ~n695 & n740 ) | ( n698 & n740 ) ;
  assign n742 = n695 | n741 ;
  assign n743 = ( x29 & n238 ) | ( x29 & n491 ) | ( n238 & n491 ) ;
  assign n744 = ~x29 & n743 ;
  assign n745 = n428 | n435 ;
  assign n746 = n49 & n419 ;
  assign n747 = n49 & n426 ;
  assign n748 = n746 | n747 ;
  assign n749 = n622 | n748 ;
  assign n750 = n49 & n499 ;
  assign n751 = ~x29 & n715 ;
  assign n752 = ( x21 & x25 ) | ( x21 & n751 ) | ( x25 & n751 ) ;
  assign n753 = ~x21 & n752 ;
  assign n754 = x30 & n753 ;
  assign n755 = n503 | n754 ;
  assign n756 = n497 | n755 ;
  assign n757 = n624 | n756 ;
  assign n758 = n750 | n757 ;
  assign n759 = n749 | n758 ;
  assign n760 = ( ~n744 & n745 ) | ( ~n744 & n759 ) | ( n745 & n759 ) ;
  assign n761 = n744 | n760 ;
  assign n762 = x3 & x20 ;
  assign n763 = ( x18 & x19 ) | ( x18 & n762 ) | ( x19 & n762 ) ;
  assign n764 = ~x18 & n763 ;
  assign n765 = x28 & n764 ;
  assign n766 = ( x21 & x22 ) | ( x21 & n765 ) | ( x22 & n765 ) ;
  assign n767 = ~x21 & n766 ;
  assign n768 = n49 & n767 ;
  assign n769 = ~x3 & x19 ;
  assign n770 = ( x2 & ~x18 ) | ( x2 & n769 ) | ( ~x18 & n769 ) ;
  assign n771 = ~x2 & n770 ;
  assign n772 = ( x21 & n260 ) | ( x21 & n771 ) | ( n260 & n771 ) ;
  assign n773 = ~x21 & n772 ;
  assign n774 = ( x29 & n111 ) | ( x29 & n773 ) | ( n111 & n773 ) ;
  assign n775 = ~x29 & n774 ;
  assign n776 = x30 & n431 ;
  assign n777 = x22 & n776 ;
  assign n778 = x23 & n776 ;
  assign n779 = n777 | n778 ;
  assign n780 = n775 | n779 ;
  assign n781 = ( ~n445 & n768 ) | ( ~n445 & n780 ) | ( n768 & n780 ) ;
  assign n782 = n445 | n781 ;
  assign n783 = n676 | n717 ;
  assign n784 = n585 | n783 ;
  assign n785 = ~x20 & n46 ;
  assign n786 = ~x21 & n785 ;
  assign n787 = ( x29 & n238 ) | ( x29 & n786 ) | ( n238 & n786 ) ;
  assign n788 = ~x29 & n787 ;
  assign n789 = x23 & ~x29 ;
  assign n790 = ( x28 & n534 ) | ( x28 & n789 ) | ( n534 & n789 ) ;
  assign n791 = ~x28 & n790 ;
  assign n792 = x30 & n791 ;
  assign n793 = ( x28 & n49 ) | ( x28 & ~n543 ) | ( n49 & ~n543 ) ;
  assign n794 = ~x28 & n793 ;
  assign n795 = n734 | n794 ;
  assign n796 = n721 | n795 ;
  assign n797 = n792 | n796 ;
  assign n798 = n788 | n797 ;
  assign n799 = x14 & ~x28 ;
  assign n800 = ( x27 & ~x29 ) | ( x27 & n799 ) | ( ~x29 & n799 ) ;
  assign n801 = ~x27 & n800 ;
  assign n802 = ~x30 & n801 ;
  assign n803 = x13 & ~x27 ;
  assign n804 = ( x14 & x21 ) | ( x14 & n803 ) | ( x21 & n803 ) ;
  assign n805 = ~x14 & n804 ;
  assign n806 = ~x29 & n805 ;
  assign n807 = ( x28 & ~x30 ) | ( x28 & n806 ) | ( ~x30 & n806 ) ;
  assign n808 = ~x28 & n807 ;
  assign n809 = n802 | n808 ;
  assign n810 = n798 | n809 ;
  assign n811 = ( ~n600 & n784 ) | ( ~n600 & n810 ) | ( n784 & n810 ) ;
  assign n812 = n600 | n811 ;
  assign n813 = x26 & ~x29 ;
  assign n814 = ( x28 & n437 ) | ( x28 & n813 ) | ( n437 & n813 ) ;
  assign n815 = ~x28 & n814 ;
  assign n816 = x30 & n815 ;
  assign n817 = ( x28 & n437 ) | ( x28 & n789 ) | ( n437 & n789 ) ;
  assign n818 = ~x28 & n817 ;
  assign n819 = x30 & n818 ;
  assign n820 = n49 & n439 ;
  assign n821 = x23 & x30 ;
  assign n822 = ( x29 & n786 ) | ( x29 & n821 ) | ( n786 & n821 ) ;
  assign n823 = ~x29 & n822 ;
  assign n824 = n452 | n823 ;
  assign n825 = n532 | n824 ;
  assign n826 = n820 | n825 ;
  assign n827 = ( ~n816 & n819 ) | ( ~n816 & n826 ) | ( n819 & n826 ) ;
  assign n828 = n816 | n827 ;
  assign n829 = n812 | n828 ;
  assign n830 = n782 | n829 ;
  assign n831 = ~x27 & n472 ;
  assign n832 = ~x28 & n831 ;
  assign n833 = n49 & n832 ;
  assign n834 = n476 | n833 ;
  assign n835 = n495 | n834 ;
  assign n836 = n469 | n835 ;
  assign n837 = n618 | n836 ;
  assign n838 = n830 | n837 ;
  assign n839 = ( ~n415 & n761 ) | ( ~n415 & n838 ) | ( n761 & n838 ) ;
  assign n840 = n415 | n839 ;
  assign n841 = x40 & ~x42 ;
  assign n842 = ( x41 & n398 ) | ( x41 & n841 ) | ( n398 & n841 ) ;
  assign n843 = ~x41 & n842 ;
  assign n844 = n388 | n843 ;
  assign n845 = n411 | n844 ;
  assign n846 = x33 & n466 ;
  assign n847 = n469 | n618 ;
  assign n848 = ( ~n458 & n846 ) | ( ~n458 & n847 ) | ( n846 & n847 ) ;
  assign n849 = n458 | n848 ;
  assign n850 = n532 | n721 ;
  assign n851 = ( ~n452 & n768 ) | ( ~n452 & n850 ) | ( n768 & n850 ) ;
  assign n852 = n452 | n851 ;
  assign n853 = n445 | n775 ;
  assign n854 = x30 & n525 ;
  assign n855 = n585 | n597 ;
  assign n856 = ( ~n636 & n638 ) | ( ~n636 & n855 ) | ( n638 & n855 ) ;
  assign n857 = n636 | n856 ;
  assign n858 = n854 | n857 ;
  assign n859 = ( n676 & ~n713 ) | ( n676 & n858 ) | ( ~n713 & n858 ) ;
  assign n860 = n713 | n859 ;
  assign n861 = n853 | n860 ;
  assign n862 = ( ~n622 & n852 ) | ( ~n622 & n861 ) | ( n852 & n861 ) ;
  assign n863 = n622 | n862 ;
  assign n864 = n497 | n745 ;
  assign n865 = n503 | n864 ;
  assign n866 = n476 | n865 ;
  assign n867 = n686 | n866 ;
  assign n868 = n863 | n867 ;
  assign n869 = ( ~n845 & n849 ) | ( ~n845 & n868 ) | ( n849 & n868 ) ;
  assign n870 = n845 | n869 ;
  assign n871 = x23 & n384 ;
  assign n872 = ( x29 & x30 ) | ( x29 & n871 ) | ( x30 & n871 ) ;
  assign n873 = ~x30 & n872 ;
  assign n874 = x31 & n873 ;
  assign n875 = ( x32 & n873 ) | ( x32 & n874 ) | ( n873 & n874 ) ;
  assign n876 = ( x29 & n384 ) | ( x29 & n821 ) | ( n384 & n821 ) ;
  assign n877 = ~x29 & n876 ;
  assign n878 = ~x32 & n873 ;
  assign n879 = ( x31 & ~x33 ) | ( x31 & n878 ) | ( ~x33 & n878 ) ;
  assign n880 = ~x31 & n879 ;
  assign n881 = x34 & n880 ;
  assign n882 = ( x35 & n880 ) | ( x35 & n881 ) | ( n880 & n881 ) ;
  assign n883 = ~x34 & n880 ;
  assign n884 = ~x35 & n883 ;
  assign n885 = ( ~x36 & n882 ) | ( ~x36 & n884 ) | ( n882 & n884 ) ;
  assign n886 = x37 & ~n885 ;
  assign n887 = ( x37 & n882 ) | ( x37 & ~n886 ) | ( n882 & ~n886 ) ;
  assign n888 = n877 | n887 ;
  assign n889 = ( ~n612 & n875 ) | ( ~n612 & n888 ) | ( n875 & n888 ) ;
  assign n890 = n612 | n889 ;
  assign n891 = x27 & x29 ;
  assign n892 = ( x28 & n472 ) | ( x28 & n891 ) | ( n472 & n891 ) ;
  assign n893 = ~x28 & n892 ;
  assign n894 = ~x30 & n893 ;
  assign n895 = ( x28 & n238 ) | ( x28 & ~n384 ) | ( n238 & ~n384 ) ;
  assign n896 = n384 & n895 ;
  assign n897 = n894 | n896 ;
  assign n898 = n133 | n480 ;
  assign n899 = ( ~x4 & x19 ) | ( ~x4 & n199 ) | ( x19 & n199 ) ;
  assign n900 = x4 & n899 ;
  assign n901 = ~x27 & x28 ;
  assign n902 = ( x21 & n900 ) | ( x21 & n901 ) | ( n900 & n901 ) ;
  assign n903 = ~x21 & n902 ;
  assign n904 = ~x30 & n903 ;
  assign n905 = x29 & n904 ;
  assign n906 = ( ~x5 & x19 ) | ( ~x5 & n199 ) | ( x19 & n199 ) ;
  assign n907 = x5 & n906 ;
  assign n908 = ~x27 & n907 ;
  assign n909 = ( x21 & ~x28 ) | ( x21 & n908 ) | ( ~x28 & n908 ) ;
  assign n910 = ~x21 & n909 ;
  assign n911 = x30 & n910 ;
  assign n912 = x29 & n911 ;
  assign n913 = n489 | n912 ;
  assign n914 = ( ~n476 & n905 ) | ( ~n476 & n913 ) | ( n905 & n913 ) ;
  assign n915 = n476 | n914 ;
  assign n916 = n898 | n915 ;
  assign n917 = ( ~n890 & n897 ) | ( ~n890 & n916 ) | ( n897 & n916 ) ;
  assign n918 = n890 | n917 ;
  assign n919 = ~x30 & n529 ;
  assign n920 = x3 & ~x18 ;
  assign n921 = ~x19 & n920 ;
  assign n922 = ~x21 & n921 ;
  assign n923 = ( x20 & ~x28 ) | ( x20 & n922 ) | ( ~x28 & n922 ) ;
  assign n924 = ~x20 & n923 ;
  assign n925 = ~x30 & n924 ;
  assign n926 = x29 & n925 ;
  assign n927 = ~x30 & n525 ;
  assign n928 = n514 | n927 ;
  assign n929 = ( ~n919 & n926 ) | ( ~n919 & n928 ) | ( n926 & n928 ) ;
  assign n930 = n919 | n929 ;
  assign n931 = n183 | n540 ;
  assign n932 = n788 | n931 ;
  assign n933 = ( x29 & n61 ) | ( x29 & n534 ) | ( n61 & n534 ) ;
  assign n934 = ~x29 & n933 ;
  assign n935 = x6 & ~x19 ;
  assign n936 = ( x3 & x18 ) | ( x3 & n935 ) | ( x18 & n935 ) ;
  assign n937 = ~x18 & n936 ;
  assign n938 = x20 & x28 ;
  assign n939 = ( x21 & n937 ) | ( x21 & n938 ) | ( n937 & n938 ) ;
  assign n940 = ~x21 & n939 ;
  assign n941 = n49 & n940 ;
  assign n942 = ~x3 & x6 ;
  assign n943 = ( x2 & ~x18 ) | ( x2 & n942 ) | ( ~x18 & n942 ) ;
  assign n944 = ~x2 & n943 ;
  assign n945 = ~x21 & n944 ;
  assign n946 = ( x19 & x20 ) | ( x19 & n945 ) | ( x20 & n945 ) ;
  assign n947 = ~x19 & n946 ;
  assign n948 = ( x29 & n111 ) | ( x29 & n947 ) | ( n111 & n947 ) ;
  assign n949 = ~x29 & n948 ;
  assign n950 = n941 | n949 ;
  assign n951 = n934 | n950 ;
  assign n952 = ( ~n537 & n932 ) | ( ~n537 & n951 ) | ( n932 & n951 ) ;
  assign n953 = n537 | n952 ;
  assign n954 = x5 & ~x18 ;
  assign n955 = ( x3 & ~x19 ) | ( x3 & n954 ) | ( ~x19 & n954 ) ;
  assign n956 = ~x3 & n955 ;
  assign n957 = ~x21 & n956 ;
  assign n958 = ( x20 & ~x28 ) | ( x20 & n957 ) | ( ~x28 & n957 ) ;
  assign n959 = ~x20 & n958 ;
  assign n960 = ~x30 & n959 ;
  assign n961 = x29 & n960 ;
  assign n962 = n549 | n961 ;
  assign n963 = ( ~n196 & n546 ) | ( ~n196 & n962 ) | ( n546 & n962 ) ;
  assign n964 = n196 | n963 ;
  assign n965 = n953 | n964 ;
  assign n966 = n930 | n965 ;
  assign n967 = ( x2 & x3 ) | ( x2 & n46 ) | ( x3 & n46 ) ;
  assign n968 = ~x3 & n967 ;
  assign n969 = ( x21 & n260 ) | ( x21 & n968 ) | ( n260 & n968 ) ;
  assign n970 = ~x21 & n969 ;
  assign n971 = ( x29 & n111 ) | ( x29 & n970 ) | ( n111 & n970 ) ;
  assign n972 = ~x29 & n971 ;
  assign n973 = n445 | n972 ;
  assign n974 = ( ~n421 & n746 ) | ( ~n421 & n973 ) | ( n746 & n973 ) ;
  assign n975 = n421 | n974 ;
  assign n976 = n501 | n865 ;
  assign n977 = ( ~n495 & n750 ) | ( ~n495 & n976 ) | ( n750 & n976 ) ;
  assign n978 = n495 | n977 ;
  assign n979 = x5 & x20 ;
  assign n980 = ( x18 & x19 ) | ( x18 & n979 ) | ( x19 & n979 ) ;
  assign n981 = ~x18 & n980 ;
  assign n982 = ~x28 & n981 ;
  assign n983 = ( x21 & x22 ) | ( x21 & n982 ) | ( x22 & n982 ) ;
  assign n984 = ~x21 & n983 ;
  assign n985 = ~x30 & n984 ;
  assign n986 = x29 & n985 ;
  assign n987 = n452 | n986 ;
  assign n988 = ( ~n441 & n532 ) | ( ~n441 & n987 ) | ( n532 & n987 ) ;
  assign n989 = n441 | n988 ;
  assign n990 = n978 | n989 ;
  assign n991 = n975 | n990 ;
  assign n992 = n568 | n585 ;
  assign n993 = n809 | n992 ;
  assign n994 = ( n594 & ~n604 ) | ( n594 & n993 ) | ( ~n604 & n993 ) ;
  assign n995 = n604 | n994 ;
  assign n996 = ( x29 & n562 ) | ( x29 & n620 ) | ( n562 & n620 ) ;
  assign n997 = ~x29 & n996 ;
  assign n998 = n107 | n997 ;
  assign n999 = ( ~n560 & n565 ) | ( ~n560 & n998 ) | ( n565 & n998 ) ;
  assign n1000 = n560 | n999 ;
  assign n1001 = n578 | n1000 ;
  assign n1002 = ( ~n676 & n995 ) | ( ~n676 & n1001 ) | ( n995 & n1001 ) ;
  assign n1003 = n676 | n1002 ;
  assign n1004 = n991 | n1003 ;
  assign n1005 = ( ~n918 & n966 ) | ( ~n918 & n1004 ) | ( n966 & n1004 ) ;
  assign n1006 = n918 | n1005 ;
  assign n1007 = n388 | n406 ;
  assign n1008 = n408 | n458 ;
  assign n1009 = n411 | n1008 ;
  assign n1010 = n133 | n682 ;
  assign n1011 = n894 | n1010 ;
  assign n1012 = n459 | n1011 ;
  assign n1013 = ( ~n469 & n477 ) | ( ~n469 & n1012 ) | ( n477 & n1012 ) ;
  assign n1014 = n469 | n1013 ;
  assign n1015 = n1009 | n1014 ;
  assign n1016 = ( ~n403 & n1007 ) | ( ~n403 & n1015 ) | ( n1007 & n1015 ) ;
  assign n1017 = n403 | n1016 ;
  assign n1018 = n744 | n864 ;
  assign n1019 = n754 | n1018 ;
  assign n1020 = ( n503 & ~n750 ) | ( n503 & n1019 ) | ( ~n750 & n1019 ) ;
  assign n1021 = n750 | n1020 ;
  assign n1022 = n775 | n972 ;
  assign n1023 = n445 | n986 ;
  assign n1024 = n768 | n1023 ;
  assign n1025 = n816 | n819 ;
  assign n1026 = n532 | n1025 ;
  assign n1027 = ( ~n452 & n1024 ) | ( ~n452 & n1026 ) | ( n1024 & n1026 ) ;
  assign n1028 = n452 | n1027 ;
  assign n1029 = n749 | n1028 ;
  assign n1030 = ( ~n777 & n1022 ) | ( ~n777 & n1029 ) | ( n1022 & n1029 ) ;
  assign n1031 = n777 | n1030 ;
  assign n1032 = n183 | n950 ;
  assign n1033 = n919 | n926 ;
  assign n1034 = n927 | n1033 ;
  assign n1035 = n593 | n1034 ;
  assign n1036 = ( ~n676 & n809 ) | ( ~n676 & n1035 ) | ( n809 & n1035 ) ;
  assign n1037 = n676 | n1036 ;
  assign n1038 = ( x29 & n238 ) | ( x29 & n534 ) | ( n238 & n534 ) ;
  assign n1039 = ~x29 & n1038 ;
  assign n1040 = x24 & n534 ;
  assign n1041 = ( x29 & x30 ) | ( x29 & n1040 ) | ( x30 & n1040 ) ;
  assign n1042 = ~x30 & n1041 ;
  assign n1043 = n961 | n1042 ;
  assign n1044 = ( ~n196 & n1039 ) | ( ~n196 & n1043 ) | ( n1039 & n1043 ) ;
  assign n1045 = n196 | n1044 ;
  assign n1046 = n1037 | n1045 ;
  assign n1047 = ( ~n1031 & n1032 ) | ( ~n1031 & n1046 ) | ( n1032 & n1046 ) ;
  assign n1048 = n1031 | n1047 ;
  assign n1049 = n905 | n913 ;
  assign n1050 = ~x30 & n832 ;
  assign n1051 = x29 & n1050 ;
  assign n1052 = n833 | n1051 ;
  assign n1053 = n686 | n1052 ;
  assign n1054 = n1049 | n1053 ;
  assign n1055 = n1048 | n1054 ;
  assign n1056 = ( ~n1017 & n1021 ) | ( ~n1017 & n1055 ) | ( n1021 & n1055 ) ;
  assign n1057 = n1017 | n1056 ;
  assign n1058 = x36 & n884 ;
  assign n1059 = ( x37 & n884 ) | ( x37 & n1058 ) | ( n884 & n1058 ) ;
  assign n1060 = n843 | n896 ;
  assign n1061 = ( ~n690 & n846 ) | ( ~n690 & n1060 ) | ( n846 & n1060 ) ;
  assign n1062 = n690 | n1061 ;
  assign n1063 = n877 | n1062 ;
  assign n1064 = ( ~n612 & n1059 ) | ( ~n612 & n1063 ) | ( n1059 & n1063 ) ;
  assign n1065 = n612 | n1064 ;
  assign n1066 = n686 | n750 ;
  assign n1067 = ( ~n501 & n503 ) | ( ~n501 & n1066 ) | ( n503 & n1066 ) ;
  assign n1068 = n501 | n1067 ;
  assign n1069 = n480 | n894 ;
  assign n1070 = n1051 | n1069 ;
  assign n1071 = ( ~n476 & n1068 ) | ( ~n476 & n1070 ) | ( n1068 & n1070 ) ;
  assign n1072 = n476 | n1071 ;
  assign n1073 = ( x29 & n111 ) | ( x29 & n562 ) | ( n111 & n562 ) ;
  assign n1074 = ~x29 & n1073 ;
  assign n1075 = n643 | n703 ;
  assign n1076 = ( ~n577 & n1074 ) | ( ~n577 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = n577 | n1076 ;
  assign n1078 = n699 | n701 ;
  assign n1079 = ( ~n854 & n1077 ) | ( ~n854 & n1078 ) | ( n1077 & n1078 ) ;
  assign n1080 = n854 | n1079 ;
  assign n1081 = ( x22 & x30 ) | ( x22 & ~n719 ) | ( x30 & ~n719 ) ;
  assign n1082 = ( n713 & n719 ) | ( n713 & n1081 ) | ( n719 & n1081 ) ;
  assign n1083 = n721 | n1082 ;
  assign n1084 = n717 | n1083 ;
  assign n1085 = n649 | n664 ;
  assign n1086 = ( ~n585 & n661 ) | ( ~n585 & n708 ) | ( n661 & n708 ) ;
  assign n1087 = n585 | n1086 ;
  assign n1088 = n559 | n638 ;
  assign n1089 = n565 | n1088 ;
  assign n1090 = n593 | n809 ;
  assign n1091 = ( ~n590 & n670 ) | ( ~n590 & n1090 ) | ( n670 & n1090 ) ;
  assign n1092 = n590 | n1091 ;
  assign n1093 = n1089 | n1092 ;
  assign n1094 = ( ~n1085 & n1087 ) | ( ~n1085 & n1093 ) | ( n1087 & n1093 ) ;
  assign n1095 = n1085 | n1094 ;
  assign n1096 = n736 | n1095 ;
  assign n1097 = ( ~n1080 & n1084 ) | ( ~n1080 & n1096 ) | ( n1084 & n1096 ) ;
  assign n1098 = n1080 | n1097 ;
  assign n1099 = n441 | n768 ;
  assign n1100 = n428 | n497 ;
  assign n1101 = ( ~n435 & n622 ) | ( ~n435 & n1100 ) | ( n622 & n1100 ) ;
  assign n1102 = n435 | n1101 ;
  assign n1103 = n746 | n779 ;
  assign n1104 = ( ~n421 & n1102 ) | ( ~n421 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = n421 | n1104 ;
  assign n1106 = n540 | n934 ;
  assign n1107 = n537 | n1106 ;
  assign n1108 = n819 | n1107 ;
  assign n1109 = n788 | n1108 ;
  assign n1110 = n1105 | n1109 ;
  assign n1111 = ( ~n853 & n1099 ) | ( ~n853 & n1110 ) | ( n1099 & n1110 ) ;
  assign n1112 = n853 | n1111 ;
  assign n1113 = n1098 | n1112 ;
  assign n1114 = ( ~n1065 & n1072 ) | ( ~n1065 & n1113 ) | ( n1072 & n1113 ) ;
  assign n1115 = n1065 | n1114 ;
  assign n1116 = n546 | n794 ;
  assign n1117 = n549 | n1116 ;
  assign n1118 = n514 | n578 ;
  assign n1119 = n1117 | n1118 ;
  assign n1120 = n792 | n934 ;
  assign n1121 = n540 | n1120 ;
  assign n1122 = ( n537 & ~n788 ) | ( n537 & n1121 ) | ( ~n788 & n1121 ) ;
  assign n1123 = n788 | n1122 ;
  assign n1124 = n560 | n568 ;
  assign n1125 = n107 | n1124 ;
  assign n1126 = n565 | n1125 ;
  assign n1127 = n1074 | n1126 ;
  assign n1128 = n590 | n604 ;
  assign n1129 = ( ~n585 & n809 ) | ( ~n585 & n1128 ) | ( n809 & n1128 ) ;
  assign n1130 = n585 | n1129 ;
  assign n1131 = n1127 | n1130 ;
  assign n1132 = ( ~n1119 & n1123 ) | ( ~n1119 & n1131 ) | ( n1123 & n1131 ) ;
  assign n1133 = n1119 | n1132 ;
  assign n1134 = x18 & ~x20 ;
  assign n1135 = ( x10 & x19 ) | ( x10 & n1134 ) | ( x19 & n1134 ) ;
  assign n1136 = ~x19 & n1135 ;
  assign n1137 = x30 & n1136 ;
  assign n1138 = ( x21 & x25 ) | ( x21 & n1137 ) | ( x25 & n1137 ) ;
  assign n1139 = ~x21 & n1138 ;
  assign n1140 = n441 | n1139 ;
  assign n1141 = n777 | n1140 ;
  assign n1142 = n421 | n1141 ;
  assign n1143 = n747 | n1142 ;
  assign n1144 = n501 | n744 ;
  assign n1145 = n754 | n1144 ;
  assign n1146 = n833 | n1145 ;
  assign n1147 = ( n480 & ~n618 ) | ( n480 & n1146 ) | ( ~n618 & n1146 ) ;
  assign n1148 = n618 | n1147 ;
  assign n1149 = ( ~x34 & x35 ) | ( ~x34 & n894 ) | ( x35 & n894 ) ;
  assign n1150 = n880 | n894 ;
  assign n1151 = ( x34 & n1149 ) | ( x34 & n1150 ) | ( n1149 & n1150 ) ;
  assign n1152 = n1059 | n1151 ;
  assign n1153 = n1148 | n1152 ;
  assign n1154 = n828 | n1153 ;
  assign n1155 = ( ~n1133 & n1143 ) | ( ~n1133 & n1154 ) | ( n1143 & n1154 ) ;
  assign n1156 = n1133 | n1155 ;
  assign n1157 = n480 | n625 ;
  assign n1158 = ( n619 & ~n833 ) | ( n619 & n1157 ) | ( ~n833 & n1157 ) ;
  assign n1159 = n833 | n1158 ;
  assign n1160 = ~x34 & x35 ;
  assign n1161 = n880 & n1160 ;
  assign n1162 = ~x32 & x33 ;
  assign n1163 = ~x31 & n873 ;
  assign n1164 = ( x32 & n1162 ) | ( x32 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1165 = n1161 | n1164 ;
  assign n1166 = n897 | n1165 ;
  assign n1167 = ( ~n612 & n1159 ) | ( ~n612 & n1166 ) | ( n1159 & n1166 ) ;
  assign n1168 = n612 | n1167 ;
  assign n1169 = n421 | n747 ;
  assign n1170 = n622 | n1169 ;
  assign n1171 = n754 | n1170 ;
  assign n1172 = ( n744 & ~n750 ) | ( n744 & n1171 ) | ( ~n750 & n1171 ) ;
  assign n1173 = n750 | n1172 ;
  assign n1174 = n537 | n792 ;
  assign n1175 = n540 | n1174 ;
  assign n1176 = n823 | n1175 ;
  assign n1177 = ( ~n452 & n788 ) | ( ~n452 & n1176 ) | ( n788 & n1176 ) ;
  assign n1178 = n452 | n1177 ;
  assign n1179 = n107 | n565 ;
  assign n1180 = n594 | n604 ;
  assign n1181 = ( ~n560 & n992 ) | ( ~n560 & n1180 ) | ( n992 & n1180 ) ;
  assign n1182 = n560 | n1181 ;
  assign n1183 = n571 | n919 ;
  assign n1184 = n927 | n1183 ;
  assign n1185 = n1182 | n1184 ;
  assign n1186 = ( ~n577 & n1179 ) | ( ~n577 & n1185 ) | ( n1179 & n1185 ) ;
  assign n1187 = n577 | n1186 ;
  assign n1188 = n549 | n1039 ;
  assign n1189 = n514 | n794 ;
  assign n1190 = n1042 | n1189 ;
  assign n1191 = ( ~n546 & n1188 ) | ( ~n546 & n1190 ) | ( n1188 & n1190 ) ;
  assign n1192 = n546 | n1191 ;
  assign n1193 = n1187 | n1192 ;
  assign n1194 = n1178 | n1193 ;
  assign n1195 = n746 | n778 ;
  assign n1196 = n775 | n1195 ;
  assign n1197 = n819 | n1196 ;
  assign n1198 = ( ~n820 & n1099 ) | ( ~n820 & n1197 ) | ( n1099 & n1197 ) ;
  assign n1199 = n820 | n1198 ;
  assign n1200 = n1194 | n1199 ;
  assign n1201 = ( ~n1168 & n1173 ) | ( ~n1168 & n1200 ) | ( n1173 & n1200 ) ;
  assign n1202 = n1168 | n1201 ;
  assign n1203 = n612 | n877 ;
  assign n1204 = n690 | n1203 ;
  assign n1205 = n403 | n843 ;
  assign n1206 = n896 | n1205 ;
  assign n1207 = ( ~n388 & n1204 ) | ( ~n388 & n1206 ) | ( n1204 & n1206 ) ;
  assign n1208 = n388 | n1207 ;
  assign n1209 = ( x31 & n873 ) | ( x31 & n1162 ) | ( n873 & n1162 ) ;
  assign n1210 = ~x31 & n1209 ;
  assign n1211 = x34 | n1210 ;
  assign n1212 = ( n880 & n1210 ) | ( n880 & n1211 ) | ( n1210 & n1211 ) ;
  assign n1213 = ( ~x36 & x37 ) | ( ~x36 & n1161 ) | ( x37 & n1161 ) ;
  assign n1214 = n884 | n1161 ;
  assign n1215 = ( x36 & n1213 ) | ( x36 & n1214 ) | ( n1213 & n1214 ) ;
  assign n1216 = n875 | n1215 ;
  assign n1217 = ( ~n1208 & n1212 ) | ( ~n1208 & n1216 ) | ( n1212 & n1216 ) ;
  assign n1218 = n1208 | n1217 ;
  assign n1219 = n469 | n846 ;
  assign n1220 = ( ~n458 & n459 ) | ( ~n458 & n1219 ) | ( n459 & n1219 ) ;
  assign n1221 = n458 | n1220 ;
  assign n1222 = n489 | n682 ;
  assign n1223 = n905 | n1222 ;
  assign n1224 = n894 | n898 ;
  assign n1225 = ( ~n477 & n1223 ) | ( ~n477 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = n477 | n1225 ;
  assign n1227 = n413 | n1226 ;
  assign n1228 = ( ~n1218 & n1221 ) | ( ~n1218 & n1227 ) | ( n1221 & n1227 ) ;
  assign n1229 = n1218 | n1228 ;
  assign n1230 = n643 | n997 ;
  assign n1231 = n577 | n1230 ;
  assign n1232 = n1074 | n1231 ;
  assign n1233 = n636 | n1232 ;
  assign n1234 = ( ~n560 & n1179 ) | ( ~n560 & n1233 ) | ( n1179 & n1233 ) ;
  assign n1235 = n560 | n1234 ;
  assign n1236 = ~x10 & n134 ;
  assign n1237 = ~x15 & n1236 ;
  assign n1238 = ( x19 & n199 ) | ( x19 & n1237 ) | ( n199 & n1237 ) ;
  assign n1239 = ~x19 & n1238 ;
  assign n1240 = x21 & n1239 ;
  assign n1241 = ( x25 & x28 ) | ( x25 & n1240 ) | ( x28 & n1240 ) ;
  assign n1242 = ~x28 & n1241 ;
  assign n1243 = n49 & n1242 ;
  assign n1244 = x5 & ~x19 ;
  assign n1245 = ( x10 & x18 ) | ( x10 & n1244 ) | ( x18 & n1244 ) ;
  assign n1246 = ~x10 & n1245 ;
  assign n1247 = ( x21 & n219 ) | ( x21 & ~n1246 ) | ( n219 & ~n1246 ) ;
  assign n1248 = n1246 & n1247 ;
  assign n1249 = ( x28 & n49 ) | ( x28 & n1248 ) | ( n49 & n1248 ) ;
  assign n1250 = ~x28 & n1249 ;
  assign n1251 = n571 | n1250 ;
  assign n1252 = ( n702 & ~n1243 ) | ( n702 & n1251 ) | ( ~n1243 & n1251 ) ;
  assign n1253 = n1243 | n1252 ;
  assign n1254 = n701 | n1253 ;
  assign n1255 = ( ~n699 & n1235 ) | ( ~n699 & n1254 ) | ( n1235 & n1254 ) ;
  assign n1256 = n699 | n1255 ;
  assign n1257 = ~x10 & x19 ;
  assign n1258 = ~x18 & n1257 ;
  assign n1259 = x21 & n1258 ;
  assign n1260 = ( x25 & x28 ) | ( x25 & n1259 ) | ( x28 & n1259 ) ;
  assign n1261 = ~x28 & n1260 ;
  assign n1262 = n49 & n1261 ;
  assign n1263 = n600 | n1262 ;
  assign n1264 = ( ~n585 & n661 ) | ( ~n585 & n1263 ) | ( n661 & n1263 ) ;
  assign n1265 = n585 | n1264 ;
  assign n1266 = ( x10 & ~x19 ) | ( x10 & n74 ) | ( ~x19 & n74 ) ;
  assign n1267 = ~x10 & n1266 ;
  assign n1268 = x25 & n1267 ;
  assign n1269 = x21 & n1268 ;
  assign n1270 = n670 | n1269 ;
  assign n1271 = n597 | n663 ;
  assign n1272 = ( n593 & ~n603 ) | ( n593 & n1271 ) | ( ~n603 & n1271 ) ;
  assign n1273 = n603 | n1272 ;
  assign n1274 = n802 | n1273 ;
  assign n1275 = ( ~n590 & n1270 ) | ( ~n590 & n1274 ) | ( n1270 & n1274 ) ;
  assign n1276 = n590 | n1275 ;
  assign n1277 = n709 | n1276 ;
  assign n1278 = ( ~n1256 & n1265 ) | ( ~n1256 & n1277 ) | ( n1265 & n1277 ) ;
  assign n1279 = n1256 | n1278 ;
  assign n1280 = ~x10 & n1135 ;
  assign n1281 = ~x29 & n1280 ;
  assign n1282 = ( x21 & x25 ) | ( x21 & n1281 ) | ( x25 & n1281 ) ;
  assign n1283 = ~x21 & n1282 ;
  assign n1284 = x30 & n1283 ;
  assign n1285 = ( x30 & n753 ) | ( x30 & n1284 ) | ( n753 & n1284 ) ;
  assign n1286 = n501 | n686 ;
  assign n1287 = n750 | n1286 ;
  assign n1288 = n912 | n1287 ;
  assign n1289 = n1052 | n1288 ;
  assign n1290 = n1018 | n1289 ;
  assign n1291 = ( ~n503 & n1285 ) | ( ~n503 & n1290 ) | ( n1285 & n1290 ) ;
  assign n1292 = n503 | n1291 ;
  assign n1293 = n816 | n1099 ;
  assign n1294 = n986 | n1293 ;
  assign n1295 = n853 | n1139 ;
  assign n1296 = ( ~n972 & n1294 ) | ( ~n972 & n1295 ) | ( n1294 & n1295 ) ;
  assign n1297 = n972 | n1296 ;
  assign n1298 = x18 & ~x19 ;
  assign n1299 = ( x10 & ~x20 ) | ( x10 & n1298 ) | ( ~x20 & n1298 ) ;
  assign n1300 = ~x10 & n1299 ;
  assign n1301 = x30 & n1300 ;
  assign n1302 = ( x21 & x25 ) | ( x21 & n1301 ) | ( x25 & n1301 ) ;
  assign n1303 = ~x21 & n1302 ;
  assign n1304 = n777 | n1303 ;
  assign n1305 = ( ~n746 & n778 ) | ( ~n746 & n1304 ) | ( n778 & n1304 ) ;
  assign n1306 = n746 | n1305 ;
  assign n1307 = n1297 | n1306 ;
  assign n1308 = ( n1170 & ~n1292 ) | ( n1170 & n1307 ) | ( ~n1292 & n1307 ) ;
  assign n1309 = n1292 | n1308 ;
  assign n1310 = ( n734 & ~n926 ) | ( n734 & n1189 ) | ( ~n926 & n1189 ) ;
  assign n1311 = n926 | n1310 ;
  assign n1312 = n961 | n1311 ;
  assign n1313 = ( ~n196 & n546 ) | ( ~n196 & n1312 ) | ( n546 & n1312 ) ;
  assign n1314 = n196 | n1313 ;
  assign n1315 = n532 | n788 ;
  assign n1316 = ( ~n183 & n823 ) | ( ~n183 & n1315 ) | ( n823 & n1315 ) ;
  assign n1317 = n183 | n1316 ;
  assign n1318 = n819 | n1317 ;
  assign n1319 = ( n452 & ~n820 ) | ( n452 & n1318 ) | ( ~n820 & n1318 ) ;
  assign n1320 = n820 | n1319 ;
  assign n1321 = ( x25 & n99 ) | ( x25 & ~n1280 ) | ( n99 & ~n1280 ) ;
  assign n1322 = n1280 & n1321 ;
  assign n1323 = ( x22 & n717 ) | ( x22 & n719 ) | ( n717 & n719 ) ;
  assign n1324 = x30 & ~n1323 ;
  assign n1325 = ( x30 & n717 ) | ( x30 & ~n1324 ) | ( n717 & ~n1324 ) ;
  assign n1326 = n721 | n1325 ;
  assign n1327 = n1322 | n1326 ;
  assign n1328 = n927 | n1327 ;
  assign n1329 = ( n529 & ~n854 ) | ( n529 & n1328 ) | ( ~n854 & n1328 ) ;
  assign n1330 = n854 | n1329 ;
  assign n1331 = n934 | n1039 ;
  assign n1332 = n792 | n1042 ;
  assign n1333 = n1331 | n1332 ;
  assign n1334 = n949 | n1333 ;
  assign n1335 = ( n537 & ~n941 ) | ( n537 & n1334 ) | ( ~n941 & n1334 ) ;
  assign n1336 = n941 | n1335 ;
  assign n1337 = n1330 | n1336 ;
  assign n1338 = ( ~n1314 & n1320 ) | ( ~n1314 & n1337 ) | ( n1320 & n1337 ) ;
  assign n1339 = n1314 | n1338 ;
  assign n1340 = n1309 | n1339 ;
  assign n1341 = ( ~n1229 & n1279 ) | ( ~n1229 & n1340 ) | ( n1279 & n1340 ) ;
  assign n1342 = n1229 | n1341 ;
  assign n1343 = n593 | n919 ;
  assign n1344 = n927 | n1343 ;
  assign n1345 = n750 | n877 ;
  assign n1346 = n833 | n1345 ;
  assign n1347 = n744 | n1346 ;
  assign n1348 = ( ~n747 & n1285 ) | ( ~n747 & n1347 ) | ( n1285 & n1347 ) ;
  assign n1349 = n747 | n1348 ;
  assign n1350 = ( x19 & ~x21 ) | ( x19 & n1134 ) | ( ~x21 & n1134 ) ;
  assign n1351 = ~x19 & n1350 ;
  assign n1352 = x30 & n1351 ;
  assign n1353 = x22 & n1352 ;
  assign n1354 = n1139 | n1353 ;
  assign n1355 = n1306 | n1354 ;
  assign n1356 = ( ~n1025 & n1349 ) | ( ~n1025 & n1355 ) | ( n1349 & n1355 ) ;
  assign n1357 = n1025 | n1356 ;
  assign n1358 = ( x29 & n534 ) | ( x29 & n595 ) | ( n534 & n595 ) ;
  assign n1359 = ~x29 & n1358 ;
  assign n1360 = n792 | n1359 ;
  assign n1361 = n1331 | n1360 ;
  assign n1362 = n823 | n1361 ;
  assign n1363 = ( n788 & ~n820 ) | ( n788 & n1362 ) | ( ~n820 & n1362 ) ;
  assign n1364 = n820 | n1363 ;
  assign n1365 = x22 & n733 ;
  assign n1366 = n794 | n1365 ;
  assign n1367 = ( ~n1243 & n1322 ) | ( ~n1243 & n1366 ) | ( n1322 & n1366 ) ;
  assign n1368 = n1243 | n1367 ;
  assign n1369 = n1262 | n1269 ;
  assign n1370 = ( n808 & ~n1250 ) | ( n808 & n1369 ) | ( ~n1250 & n1369 ) ;
  assign n1371 = n1250 | n1370 ;
  assign n1372 = n1368 | n1371 ;
  assign n1373 = ( ~n1357 & n1364 ) | ( ~n1357 & n1372 ) | ( n1364 & n1372 ) ;
  assign n1374 = n1357 | n1373 ;
  assign n1375 = n792 | n794 ;
  assign n1376 = ( ~n820 & n833 ) | ( ~n820 & n1375 ) | ( n833 & n1375 ) ;
  assign n1377 = n820 | n1376 ;
  assign n1378 = n961 | n1032 ;
  assign n1379 = ( ~n196 & n926 ) | ( ~n196 & n1378 ) | ( n926 & n1378 ) ;
  assign n1380 = n196 | n1379 ;
  assign n1381 = n912 | n986 ;
  assign n1382 = n972 | n1381 ;
  assign n1383 = n905 | n1382 ;
  assign n1384 = ( ~n133 & n1380 ) | ( ~n133 & n1383 ) | ( n1380 & n1383 ) ;
  assign n1385 = n133 | n1384 ;
  assign n1386 = n661 | n663 ;
  assign n1387 = n1262 | n1386 ;
  assign n1388 = ( x7 & x16 ) | ( x7 & n46 ) | ( x16 & n46 ) ;
  assign n1389 = ~x16 & n1388 ;
  assign n1390 = ( x21 & n260 ) | ( x21 & ~n1389 ) | ( n260 & ~n1389 ) ;
  assign n1391 = n1389 & n1390 ;
  assign n1392 = ( x29 & n620 ) | ( x29 & n1391 ) | ( n620 & n1391 ) ;
  assign n1393 = ~x29 & n1392 ;
  assign n1394 = x16 & x19 ;
  assign n1395 = ( x8 & x18 ) | ( x8 & n1394 ) | ( x18 & n1394 ) ;
  assign n1396 = ~x18 & n1395 ;
  assign n1397 = ( x21 & n260 ) | ( x21 & ~n1396 ) | ( n260 & ~n1396 ) ;
  assign n1398 = n1396 & n1397 ;
  assign n1399 = ( x29 & n620 ) | ( x29 & n1398 ) | ( n620 & n1398 ) ;
  assign n1400 = ~x29 & n1399 ;
  assign n1401 = x21 & n981 ;
  assign n1402 = ( x22 & x28 ) | ( x22 & n1401 ) | ( x28 & n1401 ) ;
  assign n1403 = ~x28 & n1402 ;
  assign n1404 = n49 & n1403 ;
  assign n1405 = n638 | n1404 ;
  assign n1406 = n655 | n1405 ;
  assign n1407 = n1400 | n1406 ;
  assign n1408 = n1393 | n1407 ;
  assign n1409 = n1387 | n1408 ;
  assign n1410 = ( ~n597 & n1270 ) | ( ~n597 & n1409 ) | ( n1270 & n1409 ) ;
  assign n1411 = n597 | n1410 ;
  assign n1412 = n690 | n896 ;
  assign n1413 = ( n873 & ~n1163 ) | ( n873 & n1412 ) | ( ~n1163 & n1412 ) ;
  assign n1414 = n721 | n1322 ;
  assign n1415 = n717 | n1414 ;
  assign n1416 = n734 | n1365 ;
  assign n1417 = n1042 | n1359 ;
  assign n1418 = n1303 | n1417 ;
  assign n1419 = ( ~n1139 & n1353 ) | ( ~n1139 & n1418 ) | ( n1353 & n1418 ) ;
  assign n1420 = n1139 | n1419 ;
  assign n1421 = n1416 | n1420 ;
  assign n1422 = ( ~n1039 & n1415 ) | ( ~n1039 & n1421 ) | ( n1415 & n1421 ) ;
  assign n1423 = n1039 | n1422 ;
  assign n1424 = n882 | n884 ;
  assign n1425 = n1164 | n1424 ;
  assign n1426 = ( ~n1413 & n1423 ) | ( ~n1413 & n1425 ) | ( n1423 & n1425 ) ;
  assign n1427 = n1413 | n1426 ;
  assign n1428 = ( x5 & x19 ) | ( x5 & n199 ) | ( x19 & n199 ) ;
  assign n1429 = ~x19 & n1428 ;
  assign n1430 = x21 & ~x28 ;
  assign n1431 = ( x25 & n1429 ) | ( x25 & n1430 ) | ( n1429 & n1430 ) ;
  assign n1432 = ~x25 & n1431 ;
  assign n1433 = n49 & n1432 ;
  assign n1434 = x5 & x10 ;
  assign n1435 = ( x18 & x19 ) | ( x18 & n1434 ) | ( x19 & n1434 ) ;
  assign n1436 = ~x19 & n1435 ;
  assign n1437 = ( x21 & n219 ) | ( x21 & ~n1436 ) | ( n219 & ~n1436 ) ;
  assign n1438 = n1436 & n1437 ;
  assign n1439 = ( x28 & n49 ) | ( x28 & n1438 ) | ( n49 & n1438 ) ;
  assign n1440 = ~x28 & n1439 ;
  assign n1441 = n1074 | n1440 ;
  assign n1442 = n1433 | n1441 ;
  assign n1443 = x7 & ~x19 ;
  assign n1444 = ( x16 & x18 ) | ( x16 & n1443 ) | ( x18 & n1443 ) ;
  assign n1445 = ~x16 & n1444 ;
  assign n1446 = ( x21 & n938 ) | ( x21 & ~n1445 ) | ( n938 & ~n1445 ) ;
  assign n1447 = n1445 & n1446 ;
  assign n1448 = x8 & x16 ;
  assign n1449 = ( x18 & x19 ) | ( x18 & n1448 ) | ( x19 & n1448 ) ;
  assign n1450 = ~x19 & n1449 ;
  assign n1451 = ( x21 & n938 ) | ( x21 & ~n1450 ) | ( n938 & ~n1450 ) ;
  assign n1452 = n1450 & n1451 ;
  assign n1453 = n1082 | n1452 ;
  assign n1454 = ( ~n699 & n1447 ) | ( ~n699 & n1453 ) | ( n1447 & n1453 ) ;
  assign n1455 = n699 | n1454 ;
  assign n1456 = n1250 | n1455 ;
  assign n1457 = ( ~n1243 & n1442 ) | ( ~n1243 & n1456 ) | ( n1442 & n1456 ) ;
  assign n1458 = n1243 | n1457 ;
  assign n1459 = n1427 | n1458 ;
  assign n1460 = n1411 | n1459 ;
  assign n1461 = n142 | n158 ;
  assign n1462 = n133 | n1461 ;
  assign n1463 = n326 | n1462 ;
  assign n1464 = ( n183 & ~n318 ) | ( n183 & n1463 ) | ( ~n318 & n1463 ) ;
  assign n1465 = n318 | n1464 ;
  assign n1466 = n257 | n296 ;
  assign n1467 = n290 | n1466 ;
  assign n1468 = ( ~n95 & n250 ) | ( ~n95 & n1467 ) | ( n250 & n1467 ) ;
  assign n1469 = n95 | n1468 ;
  assign n1470 = n113 | n264 ;
  assign n1471 = n107 | n1470 ;
  assign n1472 = n280 | n1471 ;
  assign n1473 = ( ~n223 & n1469 ) | ( ~n223 & n1472 ) | ( n1469 & n1472 ) ;
  assign n1474 = n223 | n1473 ;
  assign n1475 = n196 | n231 ;
  assign n1476 = n188 | n1475 ;
  assign n1477 = n213 | n1476 ;
  assign n1478 = ( n101 & ~n205 ) | ( n101 & n1477 ) | ( ~n205 & n1477 ) ;
  assign n1479 = n205 | n1478 ;
  assign n1480 = n1474 | n1479 ;
  assign n1481 = n1465 | n1480 ;
  assign n1482 = n305 | n312 ;
  assign n1483 = n333 | n1482 ;
  assign n1484 = n125 | n343 ;
  assign n1485 = n150 | n1484 ;
  assign n1486 = n1483 | n1485 ;
  assign n1487 = n312 | n349 ;
  assign n1488 = n356 | n1487 ;
  assign n1489 = n150 | n172 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = ~x13 & x21 ;
  assign n1492 = ( x12 & ~x14 ) | ( x12 & n1491 ) | ( ~x14 & n1491 ) ;
  assign n1493 = ~x12 & n1492 ;
  assign n1494 = ~x28 & n1493 ;
  assign n1495 = ( x27 & ~x29 ) | ( x27 & n1494 ) | ( ~x29 & n1494 ) ;
  assign n1496 = ~x27 & n1495 ;
  assign n1497 = ~x30 & n1496 ;
  assign n1498 = n898 | n905 ;
  assign n1499 = ( ~n476 & n912 ) | ( ~n476 & n1498 ) | ( n912 & n1498 ) ;
  assign n1500 = n476 | n1499 ;
  assign n1501 = n408 | n459 ;
  assign n1502 = n458 | n1501 ;
  assign n1503 = n403 | n845 ;
  assign n1504 = n612 | n1503 ;
  assign n1505 = x31 & n466 ;
  assign n1506 = ( ~x33 & n466 ) | ( ~x33 & n1505 ) | ( n466 & n1505 ) ;
  assign n1507 = n1504 | n1506 ;
  assign n1508 = n1502 | n1507 ;
  assign n1509 = n73 | n87 ;
  assign n1510 = n568 | n1509 ;
  assign n1511 = ( n113 & ~n636 ) | ( n113 & n1510 ) | ( ~n636 & n1510 ) ;
  assign n1512 = n636 | n1511 ;
  assign n1513 = n546 | n854 ;
  assign n1514 = n700 | n1513 ;
  assign n1515 = n1230 | n1514 ;
  assign n1516 = ( ~n702 & n1512 ) | ( ~n702 & n1515 ) | ( n1512 & n1515 ) ;
  assign n1517 = n702 | n1516 ;
  assign n1518 = n349 | n622 ;
  assign n1519 = n356 | n1518 ;
  assign n1520 = x30 & n488 ;
  assign n1521 = n142 | n489 ;
  assign n1522 = n171 | n1521 ;
  assign n1523 = n150 | n1522 ;
  assign n1524 = ( ~n846 & n1520 ) | ( ~n846 & n1523 ) | ( n1520 & n1523 ) ;
  assign n1525 = n846 | n1524 ;
  assign n1526 = n625 | n1525 ;
  assign n1527 = ( ~n165 & n1519 ) | ( ~n165 & n1526 ) | ( n1519 & n1526 ) ;
  assign n1528 = n165 | n1527 ;
  assign n1529 = ( x29 & n534 ) | ( x29 & n620 ) | ( n534 & n620 ) ;
  assign n1530 = ~x29 & n1529 ;
  assign n1531 = ( x29 & ~n543 ) | ( x29 & n620 ) | ( ~n543 & n620 ) ;
  assign n1532 = ~x29 & n1531 ;
  assign n1533 = n196 | n1532 ;
  assign n1534 = n537 | n1533 ;
  assign n1535 = n183 | n1534 ;
  assign n1536 = ( ~n441 & n1530 ) | ( ~n441 & n1535 ) | ( n1530 & n1535 ) ;
  assign n1537 = n441 | n1536 ;
  assign n1538 = ~x29 & n443 ;
  assign n1539 = ~x30 & n1538 ;
  assign n1540 = n768 | n1539 ;
  assign n1541 = n312 | n1540 ;
  assign n1542 = n775 | n1541 ;
  assign n1543 = ( ~n421 & n1537 ) | ( ~n421 & n1542 ) | ( n1537 & n1542 ) ;
  assign n1544 = n421 | n1543 ;
  assign n1545 = n1528 | n1544 ;
  assign n1546 = ( ~n1508 & n1517 ) | ( ~n1508 & n1545 ) | ( n1517 & n1545 ) ;
  assign n1547 = n1508 | n1546 ;
  assign n1548 = x3 | x18 ;
  assign n1549 = ( ~x2 & x6 ) | ( ~x2 & n1548 ) | ( x6 & n1548 ) ;
  assign n1550 = x2 | n1549 ;
  assign n1551 = x21 | n1550 ;
  assign n1552 = ( x19 & x20 ) | ( x19 & ~n1551 ) | ( x20 & ~n1551 ) ;
  assign n1553 = ~x19 & n1552 ;
  assign n1554 = ( x29 & n111 ) | ( x29 & n1553 ) | ( n111 & n1553 ) ;
  assign n1555 = ~x29 & n1554 ;
  assign n1556 = n183 | n1555 ;
  assign n1557 = n788 | n1556 ;
  assign n1558 = n445 | n768 ;
  assign n1559 = ( n312 & ~n318 ) | ( n312 & n1558 ) | ( ~n318 & n1558 ) ;
  assign n1560 = n318 | n1559 ;
  assign n1561 = n823 | n1560 ;
  assign n1562 = ( ~n820 & n1557 ) | ( ~n820 & n1561 ) | ( n1557 & n1561 ) ;
  assign n1563 = n820 | n1562 ;
  assign n1564 = n334 | n775 ;
  assign n1565 = ( ~n746 & n747 ) | ( ~n746 & n1564 ) | ( n747 & n1564 ) ;
  assign n1566 = n746 | n1565 ;
  assign n1567 = n305 | n744 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = ( n357 & ~n1563 ) | ( n357 & n1568 ) | ( ~n1563 & n1568 ) ;
  assign n1570 = n1563 | n1569 ;
  assign n1571 = n158 | n750 ;
  assign n1572 = n343 | n1571 ;
  assign n1573 = ( ~n125 & n754 ) | ( ~n125 & n1572 ) | ( n754 & n1572 ) ;
  assign n1574 = n125 | n1573 ;
  assign n1575 = n1052 | n1574 ;
  assign n1576 = n172 | n1575 ;
  assign n1577 = n477 | n877 ;
  assign n1578 = ( ~n406 & n480 ) | ( ~n406 & n1577 ) | ( n480 & n1577 ) ;
  assign n1579 = n406 | n1578 ;
  assign n1580 = n905 | n1520 ;
  assign n1581 = n912 | n1580 ;
  assign n1582 = n150 | n1581 ;
  assign n1583 = n618 | n1582 ;
  assign n1584 = n1579 | n1583 ;
  assign n1585 = ( ~n1570 & n1576 ) | ( ~n1570 & n1584 ) | ( n1576 & n1584 ) ;
  assign n1586 = n1570 | n1585 ;
  assign n1587 = n240 | n590 ;
  assign n1588 = n257 | n604 ;
  assign n1589 = ( ~n95 & n593 ) | ( ~n95 & n1588 ) | ( n593 & n1588 ) ;
  assign n1590 = n95 | n1589 ;
  assign n1591 = n297 | n1590 ;
  assign n1592 = ( ~n249 & n1587 ) | ( ~n249 & n1591 ) | ( n1587 & n1591 ) ;
  assign n1593 = n249 | n1592 ;
  assign n1594 = n279 | n577 ;
  assign n1595 = n264 | n560 ;
  assign n1596 = n568 | n1595 ;
  assign n1597 = ( n113 & ~n585 ) | ( n113 & n1596 ) | ( ~n585 & n1596 ) ;
  assign n1598 = n585 | n1597 ;
  assign n1599 = n1179 | n1598 ;
  assign n1600 = ( ~n1593 & n1594 ) | ( ~n1593 & n1599 ) | ( n1594 & n1599 ) ;
  assign n1601 = n1593 | n1600 ;
  assign n1602 = n101 | n919 ;
  assign n1603 = ( ~n205 & n927 ) | ( ~n205 & n1602 ) | ( n927 & n1602 ) ;
  assign n1604 = n205 | n1603 ;
  assign n1605 = n223 | n571 ;
  assign n1606 = n272 | n1605 ;
  assign n1607 = n676 | n1606 ;
  assign n1608 = ( ~n213 & n1604 ) | ( ~n213 & n1607 ) | ( n1604 & n1607 ) ;
  assign n1609 = n213 | n1608 ;
  assign n1610 = ( x6 & ~x19 ) | ( x6 & n920 ) | ( ~x19 & n920 ) ;
  assign n1611 = ~x6 & n1610 ;
  assign n1612 = ( x21 & n938 ) | ( x21 & n1611 ) | ( n938 & n1611 ) ;
  assign n1613 = ~x21 & n1612 ;
  assign n1614 = n49 & n1613 ;
  assign n1615 = x3 | x19 ;
  assign n1616 = ( ~x2 & x18 ) | ( ~x2 & n1615 ) | ( x18 & n1615 ) ;
  assign n1617 = x2 | n1616 ;
  assign n1618 = x20 | n1617 ;
  assign n1619 = x21 | n1618 ;
  assign n1620 = ( x29 & n111 ) | ( x29 & ~n1619 ) | ( n111 & ~n1619 ) ;
  assign n1621 = ~x29 & n1620 ;
  assign n1622 = n231 | n1189 ;
  assign n1623 = ( ~n196 & n1621 ) | ( ~n196 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = n196 | n1623 ;
  assign n1625 = n1614 | n1624 ;
  assign n1626 = ( ~n188 & n1120 ) | ( ~n188 & n1625 ) | ( n1120 & n1625 ) ;
  assign n1627 = n188 | n1626 ;
  assign n1628 = n1609 | n1627 ;
  assign n1629 = ( ~n1586 & n1601 ) | ( ~n1586 & n1628 ) | ( n1601 & n1628 ) ;
  assign n1630 = n1586 | n1629 ;
  assign n1631 = n489 | n1051 ;
  assign n1632 = n624 | n1631 ;
  assign n1633 = n133 | n618 ;
  assign n1634 = n150 | n1633 ;
  assign n1635 = n406 | n1634 ;
  assign n1636 = ( ~n843 & n846 ) | ( ~n843 & n1635 ) | ( n846 & n1635 ) ;
  assign n1637 = n843 | n1636 ;
  assign n1638 = n1484 | n1637 ;
  assign n1639 = ( ~n158 & n1632 ) | ( ~n158 & n1638 ) | ( n1632 & n1638 ) ;
  assign n1640 = n158 | n1639 ;
  assign n1641 = ( x14 & ~x20 ) | ( x14 & n1298 ) | ( ~x20 & n1298 ) ;
  assign n1642 = ~x14 & n1641 ;
  assign n1643 = ~x27 & n1642 ;
  assign n1644 = ( x21 & ~x28 ) | ( x21 & n1643 ) | ( ~x28 & n1643 ) ;
  assign n1645 = ~x21 & n1644 ;
  assign n1646 = ~x29 & n1645 ;
  assign n1647 = ~x30 & n1646 ;
  assign n1648 = ( x14 & ~x19 ) | ( x14 & n74 ) | ( ~x19 & n74 ) ;
  assign n1649 = ~x14 & n1648 ;
  assign n1650 = ~x23 & n1649 ;
  assign n1651 = ( x21 & ~x27 ) | ( x21 & n1650 ) | ( ~x27 & n1650 ) ;
  assign n1652 = ~x21 & n1651 ;
  assign n1653 = ~x29 & n1652 ;
  assign n1654 = ( x28 & ~x30 ) | ( x28 & n1653 ) | ( ~x30 & n1653 ) ;
  assign n1655 = ~x28 & n1654 ;
  assign n1656 = x13 & ~x21 ;
  assign n1657 = ( x14 & ~x27 ) | ( x14 & n1656 ) | ( ~x27 & n1656 ) ;
  assign n1658 = ~x14 & n1657 ;
  assign n1659 = ~x29 & n1658 ;
  assign n1660 = ( x28 & ~x30 ) | ( x28 & n1659 ) | ( ~x30 & n1659 ) ;
  assign n1661 = ~x28 & n1660 ;
  assign n1662 = n1655 | n1661 ;
  assign n1663 = ( ~n1497 & n1647 ) | ( ~n1497 & n1662 ) | ( n1647 & n1662 ) ;
  assign n1664 = n1497 | n1663 ;
  assign n1665 = ( x5 & x15 ) | ( x5 & n46 ) | ( x15 & n46 ) ;
  assign n1666 = ~x5 & n1665 ;
  assign n1667 = ( x21 & n260 ) | ( x21 & ~n1666 ) | ( n260 & ~n1666 ) ;
  assign n1668 = n1666 & n1667 ;
  assign n1669 = ( x28 & n49 ) | ( x28 & n1668 ) | ( n49 & n1668 ) ;
  assign n1670 = ~x28 & n1669 ;
  assign n1671 = ( ~n560 & n1510 ) | ( ~n560 & n1670 ) | ( n1510 & n1670 ) ;
  assign n1672 = n560 | n1671 ;
  assign n1673 = n1664 | n1672 ;
  assign n1674 = ( n594 & ~n603 ) | ( n594 & n1673 ) | ( ~n603 & n1673 ) ;
  assign n1675 = n603 | n1674 ;
  assign n1676 = n333 | n622 ;
  assign n1677 = n312 | n1539 ;
  assign n1678 = n326 | n1677 ;
  assign n1679 = n231 | n1532 ;
  assign n1680 = ( n514 & ~n919 ) | ( n514 & n1679 ) | ( ~n919 & n1679 ) ;
  assign n1681 = n919 | n1680 ;
  assign n1682 = n188 | n1681 ;
  assign n1683 = ( ~n318 & n1530 ) | ( ~n318 & n1682 ) | ( n1530 & n1682 ) ;
  assign n1684 = n318 | n1683 ;
  assign n1685 = n1678 | n1684 ;
  assign n1686 = ( ~n305 & n1676 ) | ( ~n305 & n1685 ) | ( n1676 & n1685 ) ;
  assign n1687 = n305 | n1686 ;
  assign n1688 = x15 & ~x19 ;
  assign n1689 = ( x5 & x18 ) | ( x5 & n1688 ) | ( x18 & n1688 ) ;
  assign n1690 = ~x5 & n1689 ;
  assign n1691 = x20 & n1690 ;
  assign n1692 = ( x21 & x28 ) | ( x21 & n1691 ) | ( x28 & n1691 ) ;
  assign n1693 = ~x28 & n1692 ;
  assign n1694 = n49 & n1693 ;
  assign n1695 = ~x16 & x19 ;
  assign n1696 = ( x7 & ~x18 ) | ( x7 & n1695 ) | ( ~x18 & n1695 ) ;
  assign n1697 = ~x7 & n1696 ;
  assign n1698 = ( x21 & n260 ) | ( x21 & ~n1697 ) | ( n260 & ~n1697 ) ;
  assign n1699 = n1697 & n1698 ;
  assign n1700 = ( x29 & n620 ) | ( x29 & n1699 ) | ( n620 & n1699 ) ;
  assign n1701 = ~x29 & n1700 ;
  assign n1702 = ( x8 & x16 ) | ( x8 & n46 ) | ( x16 & n46 ) ;
  assign n1703 = ~x8 & n1702 ;
  assign n1704 = ( x21 & n260 ) | ( x21 & ~n1703 ) | ( n260 & ~n1703 ) ;
  assign n1705 = n1703 & n1704 ;
  assign n1706 = ( x29 & n620 ) | ( x29 & n1705 ) | ( n620 & n1705 ) ;
  assign n1707 = ~x29 & n1706 ;
  assign n1708 = n565 | n1707 ;
  assign n1709 = n1701 | n1708 ;
  assign n1710 = n1694 | n1709 ;
  assign n1711 = ( ~n577 & n997 ) | ( ~n577 & n1710 ) | ( n997 & n1710 ) ;
  assign n1712 = n577 | n1711 ;
  assign n1713 = ~x16 & x18 ;
  assign n1714 = ( x7 & ~x19 ) | ( x7 & n1713 ) | ( ~x19 & n1713 ) ;
  assign n1715 = ~x7 & n1714 ;
  assign n1716 = ( x21 & n938 ) | ( x21 & ~n1715 ) | ( n938 & ~n1715 ) ;
  assign n1717 = n1715 & n1716 ;
  assign n1718 = x16 & ~x19 ;
  assign n1719 = ( x8 & x18 ) | ( x8 & n1718 ) | ( x18 & n1718 ) ;
  assign n1720 = ~x8 & n1719 ;
  assign n1721 = ( x21 & n938 ) | ( x21 & ~n1720 ) | ( n938 & ~n1720 ) ;
  assign n1722 = n1720 & n1721 ;
  assign n1723 = n571 | n1722 ;
  assign n1724 = n1717 | n1723 ;
  assign n1725 = n701 | n1724 ;
  assign n1726 = ( ~n927 & n1712 ) | ( ~n927 & n1725 ) | ( n1712 & n1725 ) ;
  assign n1727 = n927 | n1726 ;
  assign n1728 = n1687 | n1727 ;
  assign n1729 = ( ~n1640 & n1675 ) | ( ~n1640 & n1728 ) | ( n1675 & n1728 ) ;
  assign n1730 = n1640 | n1729 ;
  assign n1731 = n1204 | n1424 ;
  assign n1732 = ( n875 & ~n1210 ) | ( n875 & n1731 ) | ( ~n1210 & n1731 ) ;
  assign n1733 = n1210 | n1732 ;
  assign n1734 = n150 | n1520 ;
  assign n1735 = n905 | n1734 ;
  assign n1736 = ( x33 & n466 ) | ( x33 & n1505 ) | ( n466 & n1505 ) ;
  assign n1737 = n477 | n1069 ;
  assign n1738 = n1736 | n1737 ;
  assign n1739 = n682 | n1738 ;
  assign n1740 = ( ~n133 & n1735 ) | ( ~n133 & n1739 ) | ( n1735 & n1739 ) ;
  assign n1741 = n133 | n1740 ;
  assign n1742 = ~x31 & n466 ;
  assign n1743 = ~x33 & n1742 ;
  assign n1744 = n459 | n1743 ;
  assign n1745 = n1009 | n1744 ;
  assign n1746 = n1205 | n1745 ;
  assign n1747 = ( ~n896 & n1007 ) | ( ~n896 & n1746 ) | ( n1007 & n1746 ) ;
  assign n1748 = n896 | n1747 ;
  assign n1749 = n165 | n624 ;
  assign n1750 = n171 | n1749 ;
  assign n1751 = n495 | n1051 ;
  assign n1752 = n833 | n1751 ;
  assign n1753 = n489 | n1752 ;
  assign n1754 = ( ~n142 & n912 ) | ( ~n142 & n1753 ) | ( n912 & n1753 ) ;
  assign n1755 = n142 | n1754 ;
  assign n1756 = n1571 | n1755 ;
  assign n1757 = ( ~n501 & n1750 ) | ( ~n501 & n1756 ) | ( n1750 & n1756 ) ;
  assign n1758 = n501 | n1757 ;
  assign n1759 = n1748 | n1758 ;
  assign n1760 = ( ~n1733 & n1741 ) | ( ~n1733 & n1759 ) | ( n1741 & n1759 ) ;
  assign n1761 = n1733 | n1760 ;
  assign n1762 = n1032 | n1614 ;
  assign n1763 = ( n1530 & ~n1555 ) | ( n1530 & n1762 ) | ( ~n1555 & n1762 ) ;
  assign n1764 = n1555 | n1763 ;
  assign n1765 = n318 | n1539 ;
  assign n1766 = n441 | n1765 ;
  assign n1767 = n312 | n1022 ;
  assign n1768 = ( ~n445 & n768 ) | ( ~n445 & n1767 ) | ( n768 & n1767 ) ;
  assign n1769 = n445 | n1768 ;
  assign n1770 = n1025 | n1769 ;
  assign n1771 = ( ~n986 & n1766 ) | ( ~n986 & n1770 ) | ( n1766 & n1770 ) ;
  assign n1772 = n986 | n1771 ;
  assign n1773 = n532 | n540 ;
  assign n1774 = n788 | n1773 ;
  assign n1775 = n452 | n1774 ;
  assign n1776 = ( ~n820 & n823 ) | ( ~n820 & n1775 ) | ( n823 & n1775 ) ;
  assign n1777 = n820 | n1776 ;
  assign n1778 = n1772 | n1777 ;
  assign n1779 = n1764 | n1778 ;
  assign n1780 = n497 | n1567 ;
  assign n1781 = ( n357 & ~n435 ) | ( n357 & n1780 ) | ( ~n435 & n1780 ) ;
  assign n1782 = n435 | n1781 ;
  assign n1783 = n779 | n1303 ;
  assign n1784 = ( ~n746 & n1354 ) | ( ~n746 & n1783 ) | ( n1354 & n1783 ) ;
  assign n1785 = n746 | n1784 ;
  assign n1786 = n326 | n1169 ;
  assign n1787 = n1785 | n1786 ;
  assign n1788 = ( ~n428 & n1676 ) | ( ~n428 & n1787 ) | ( n1676 & n1787 ) ;
  assign n1789 = n428 | n1788 ;
  assign n1790 = n343 | n1285 ;
  assign n1791 = ( ~n125 & n503 ) | ( ~n125 & n1790 ) | ( n503 & n1790 ) ;
  assign n1792 = n125 | n1791 ;
  assign n1793 = n1789 | n1792 ;
  assign n1794 = ( ~n1779 & n1782 ) | ( ~n1779 & n1793 ) | ( n1782 & n1793 ) ;
  assign n1795 = n1779 | n1794 ;
  assign n1796 = n213 | n699 ;
  assign n1797 = n927 | n1796 ;
  assign n1798 = n676 | n1797 ;
  assign n1799 = ( ~n223 & n700 ) | ( ~n223 & n1798 ) | ( n700 & n1798 ) ;
  assign n1800 = n223 | n1799 ;
  assign n1801 = n919 | n1082 ;
  assign n1802 = ( ~n205 & n854 ) | ( ~n205 & n1801 ) | ( n854 & n1801 ) ;
  assign n1803 = n205 | n1802 ;
  assign n1804 = n272 | n1722 ;
  assign n1805 = n571 | n1804 ;
  assign n1806 = n1452 | n1805 ;
  assign n1807 = ( ~n1243 & n1447 ) | ( ~n1243 & n1806 ) | ( n1447 & n1806 ) ;
  assign n1808 = n1243 | n1807 ;
  assign n1809 = n702 | n1717 ;
  assign n1810 = n1694 | n1809 ;
  assign n1811 = n1440 | n1810 ;
  assign n1812 = ( ~n1250 & n1433 ) | ( ~n1250 & n1811 ) | ( n1433 & n1811 ) ;
  assign n1813 = n1250 | n1812 ;
  assign n1814 = n1808 | n1813 ;
  assign n1815 = ( ~n1800 & n1803 ) | ( ~n1800 & n1814 ) | ( n1803 & n1814 ) ;
  assign n1816 = n1800 | n1815 ;
  assign n1817 = n794 | n926 ;
  assign n1818 = n734 | n1817 ;
  assign n1819 = n961 | n1818 ;
  assign n1820 = ( ~n231 & n546 ) | ( ~n231 & n1819 ) | ( n546 & n1819 ) ;
  assign n1821 = n231 | n1820 ;
  assign n1822 = n1533 | n1621 ;
  assign n1823 = n792 | n1417 ;
  assign n1824 = ( ~n188 & n537 ) | ( ~n188 & n1823 ) | ( n537 & n1823 ) ;
  assign n1825 = n188 | n1824 ;
  assign n1826 = n1822 | n1825 ;
  assign n1827 = ( ~n934 & n1188 ) | ( ~n934 & n1826 ) | ( n1188 & n1826 ) ;
  assign n1828 = n934 | n1827 ;
  assign n1829 = n514 | n1415 ;
  assign n1830 = ( ~n101 & n1365 ) | ( ~n101 & n1829 ) | ( n1365 & n1829 ) ;
  assign n1831 = n101 | n1830 ;
  assign n1832 = n1828 | n1831 ;
  assign n1833 = ( ~n1816 & n1821 ) | ( ~n1816 & n1832 ) | ( n1821 & n1832 ) ;
  assign n1834 = n1816 | n1833 ;
  assign n1835 = n1179 | n1393 ;
  assign n1836 = n1707 | n1835 ;
  assign n1837 = ( ~n1400 & n1701 ) | ( ~n1400 & n1836 ) | ( n1701 & n1836 ) ;
  assign n1838 = n1400 | n1837 ;
  assign n1839 = n1594 | n1838 ;
  assign n1840 = ( ~n1074 & n1230 ) | ( ~n1074 & n1839 ) | ( n1230 & n1839 ) ;
  assign n1841 = n1074 | n1840 ;
  assign n1842 = n73 | n663 ;
  assign n1843 = n70 | n1842 ;
  assign n1844 = n95 | n597 ;
  assign n1845 = n603 | n1844 ;
  assign n1846 = n593 | n1466 ;
  assign n1847 = n1845 | n1846 ;
  assign n1848 = n600 | n1847 ;
  assign n1849 = ( ~n51 & n1843 ) | ( ~n51 & n1848 ) | ( n1843 & n1848 ) ;
  assign n1850 = n51 | n1849 ;
  assign n1851 = n585 | n1262 ;
  assign n1852 = n661 | n1851 ;
  assign n1853 = n655 | n1852 ;
  assign n1854 = ( n113 & ~n568 ) | ( n113 & n1853 ) | ( ~n568 & n1853 ) ;
  assign n1855 = n568 | n1854 ;
  assign n1856 = n638 | n1670 ;
  assign n1857 = n1404 | n1856 ;
  assign n1858 = n1855 | n1857 ;
  assign n1859 = ( ~n636 & n1595 ) | ( ~n636 & n1858 ) | ( n1595 & n1858 ) ;
  assign n1860 = n636 | n1859 ;
  assign n1861 = n249 | n1269 ;
  assign n1862 = n290 | n1861 ;
  assign n1863 = x26 & n99 ;
  assign n1864 = ( x19 & n199 ) | ( x19 & ~n1863 ) | ( n199 & ~n1863 ) ;
  assign n1865 = n1863 & n1864 ;
  assign n1866 = n1655 | n1865 ;
  assign n1867 = n802 | n1866 ;
  assign n1868 = n1647 | n1867 ;
  assign n1869 = ( ~n1497 & n1661 ) | ( ~n1497 & n1868 ) | ( n1661 & n1868 ) ;
  assign n1870 = n1497 | n1869 ;
  assign n1871 = n1587 | n1870 ;
  assign n1872 = ( ~n670 & n1862 ) | ( ~n670 & n1871 ) | ( n1862 & n1871 ) ;
  assign n1873 = n670 | n1872 ;
  assign n1874 = n1860 | n1873 ;
  assign n1875 = ( ~n1841 & n1850 ) | ( ~n1841 & n1874 ) | ( n1850 & n1874 ) ;
  assign n1876 = n1841 | n1875 ;
  assign n1877 = n1834 | n1876 ;
  assign n1878 = ( ~n1761 & n1795 ) | ( ~n1761 & n1877 ) | ( n1795 & n1877 ) ;
  assign n1879 = n1761 | n1878 ;
  assign n1880 = x21 & n49 ;
  assign n1881 = ( x18 & n90 ) | ( x18 & n1880 ) | ( n90 & n1880 ) ;
  assign n1882 = ~x18 & n1881 ;
  assign n1883 = ~x21 & x29 ;
  assign n1884 = ~x30 & n1883 ;
  assign n1885 = x18 & n1884 ;
  assign n1886 = ( x19 & x20 ) | ( x19 & n1885 ) | ( x20 & n1885 ) ;
  assign n1887 = ~x20 & n1886 ;
  assign n1888 = n1882 | n1887 ;
  assign n1889 = x25 & n1888 ;
  assign n1890 = ( x22 & n1888 ) | ( x22 & n1889 ) | ( n1888 & n1889 ) ;
  assign n1891 = ~x19 & x28 ;
  assign n1892 = x11 & x30 ;
  assign n1893 = ( x26 & ~n1891 ) | ( x26 & n1892 ) | ( ~n1891 & n1892 ) ;
  assign n1894 = n1891 & n1893 ;
  assign n1895 = ( x3 & x19 ) | ( x3 & n1894 ) | ( x19 & n1894 ) ;
  assign n1896 = x27 & ~n1895 ;
  assign n1897 = ( x27 & n1894 ) | ( x27 & ~n1896 ) | ( n1894 & ~n1896 ) ;
  assign n1898 = x18 & ~n1897 ;
  assign n1899 = ~x3 & x30 ;
  assign n1900 = x2 & n1899 ;
  assign n1901 = n1891 & n1900 ;
  assign n1902 = x18 | n1901 ;
  assign n1903 = ~n1898 & n1902 ;
  assign n1904 = ~x29 & n1903 ;
  assign n1905 = x22 & x28 ;
  assign n1906 = ( ~x5 & x22 ) | ( ~x5 & n1905 ) | ( x22 & n1905 ) ;
  assign n1907 = x19 & ~n1906 ;
  assign n1908 = x23 & ~x28 ;
  assign n1909 = x19 | n1908 ;
  assign n1910 = ~n1907 & n1909 ;
  assign n1911 = ( x18 & ~x30 ) | ( x18 & n1910 ) | ( ~x30 & n1910 ) ;
  assign n1912 = x4 | x27 ;
  assign n1913 = x19 & ~x28 ;
  assign n1914 = x19 & ~n1913 ;
  assign n1915 = ~n1912 & n1914 ;
  assign n1916 = ( x26 & ~n1913 ) | ( x26 & n1914 ) | ( ~n1913 & n1914 ) ;
  assign n1917 = ( ~x28 & n1915 ) | ( ~x28 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = ( x18 & x30 ) | ( x18 & ~n1917 ) | ( x30 & ~n1917 ) ;
  assign n1919 = n1911 & ~n1918 ;
  assign n1920 = ~x5 & x30 ;
  assign n1921 = ~x27 & n1920 ;
  assign n1922 = x18 & n1921 ;
  assign n1923 = ( x19 & x28 ) | ( x19 & n1922 ) | ( x28 & n1922 ) ;
  assign n1924 = ~x28 & n1923 ;
  assign n1925 = n1919 | n1924 ;
  assign n1926 = x29 & n1925 ;
  assign n1927 = n1904 | n1926 ;
  assign n1928 = x20 & n1927 ;
  assign n1929 = ( ~x26 & x28 ) | ( ~x26 & x29 ) | ( x28 & x29 ) ;
  assign n1930 = ( x29 & x30 ) | ( x29 & ~n1929 ) | ( x30 & ~n1929 ) ;
  assign n1931 = ( ~x28 & x30 ) | ( ~x28 & n1929 ) | ( x30 & n1929 ) ;
  assign n1932 = n1930 & ~n1931 ;
  assign n1933 = x19 & ~n46 ;
  assign n1934 = n1932 & n1933 ;
  assign n1935 = ~x28 & x29 ;
  assign n1936 = ( x5 & ~x30 ) | ( x5 & n1935 ) | ( ~x30 & n1935 ) ;
  assign n1937 = ~x5 & n1936 ;
  assign n1938 = ( x2 & x28 ) | ( x2 & n49 ) | ( x28 & n49 ) ;
  assign n1939 = ~x2 & n1938 ;
  assign n1940 = ~x3 & n1939 ;
  assign n1941 = ( ~x3 & n1937 ) | ( ~x3 & n1940 ) | ( n1937 & n1940 ) ;
  assign n1942 = ( ~n46 & n1933 ) | ( ~n46 & n1941 ) | ( n1933 & n1941 ) ;
  assign n1943 = ( ~x18 & n1934 ) | ( ~x18 & n1942 ) | ( n1934 & n1942 ) ;
  assign n1944 = x20 | n1943 ;
  assign n1945 = ( ~x20 & n1928 ) | ( ~x20 & n1944 ) | ( n1928 & n1944 ) ;
  assign n1946 = x21 | n1945 ;
  assign n1947 = x5 | x28 ;
  assign n1948 = x15 | n1947 ;
  assign n1949 = ( x20 & x22 ) | ( x20 & x28 ) | ( x22 & x28 ) ;
  assign n1950 = n1948 | n1949 ;
  assign n1951 = ( x28 & ~n1948 ) | ( x28 & n1950 ) | ( ~n1948 & n1950 ) ;
  assign n1952 = x19 & ~n1951 ;
  assign n1953 = x19 | n254 ;
  assign n1954 = ~n1952 & n1953 ;
  assign n1955 = ( x18 & ~x30 ) | ( x18 & n1954 ) | ( ~x30 & n1954 ) ;
  assign n1956 = ( x19 & n199 ) | ( x19 & ~n1948 ) | ( n199 & ~n1948 ) ;
  assign n1957 = ~x19 & n1956 ;
  assign n1958 = x30 & n1957 ;
  assign n1959 = ( n1954 & ~n1955 ) | ( n1954 & n1958 ) | ( ~n1955 & n1958 ) ;
  assign n1960 = ~x29 & n1959 ;
  assign n1961 = x21 & ~n1960 ;
  assign n1962 = n1946 & ~n1961 ;
  assign n1963 = ~x22 & x23 ;
  assign n1964 = x28 | x29 ;
  assign n1965 = x30 & n1964 ;
  assign n1966 = ( n99 & n1883 ) | ( n99 & ~n1965 ) | ( n1883 & ~n1965 ) ;
  assign n1967 = ~x20 & n1966 ;
  assign n1968 = ( x22 & n1963 ) | ( x22 & n1967 ) | ( n1963 & n1967 ) ;
  assign n1969 = ( x1 & n46 ) | ( x1 & n1968 ) | ( n46 & n1968 ) ;
  assign n1970 = ~x1 & n1969 ;
  assign n1971 = n57 | n1970 ;
  assign n1972 = ( ~n63 & n80 ) | ( ~n63 & n1971 ) | ( n80 & n1971 ) ;
  assign n1973 = n63 | n1972 ;
  assign n1974 = ( ~n1890 & n1962 ) | ( ~n1890 & n1973 ) | ( n1962 & n1973 ) ;
  assign n1975 = x0 & ~n1973 ;
  assign n1976 = ( n1890 & n1974 ) | ( n1890 & ~n1975 ) | ( n1974 & ~n1975 ) ;
  assign n1977 = n865 | n905 ;
  assign n1978 = ( n480 & ~n495 ) | ( n480 & n1977 ) | ( ~n495 & n1977 ) ;
  assign n1979 = n495 | n1978 ;
  assign n1980 = n565 | n571 ;
  assign n1981 = ( n577 & ~n676 ) | ( n577 & n1980 ) | ( ~n676 & n1980 ) ;
  assign n1982 = n676 | n1981 ;
  assign n1983 = n927 | n1982 ;
  assign n1984 = ( n514 & ~n919 ) | ( n514 & n1983 ) | ( ~n919 & n1983 ) ;
  assign n1985 = n919 | n1984 ;
  assign n1986 = n540 | n549 ;
  assign n1987 = ( ~n532 & n537 ) | ( ~n532 & n1986 ) | ( n537 & n1986 ) ;
  assign n1988 = n532 | n1987 ;
  assign n1989 = n972 | n1988 ;
  assign n1990 = ( ~n452 & n986 ) | ( ~n452 & n1989 ) | ( n986 & n1989 ) ;
  assign n1991 = n452 | n1990 ;
  assign n1992 = n1985 | n1991 ;
  assign n1993 = ( n1182 & ~n1979 ) | ( n1182 & n1992 ) | ( ~n1979 & n1992 ) ;
  assign n1994 = n1979 | n1993 ;
  assign n1995 = n1404 | n1433 ;
  assign n1996 = ( ~n926 & n1440 ) | ( ~n926 & n1995 ) | ( n1440 & n1995 ) ;
  assign n1997 = n926 | n1996 ;
  assign n1998 = n912 | n1997 ;
  assign n1999 = ( ~n961 & n986 ) | ( ~n961 & n1998 ) | ( n986 & n1998 ) ;
  assign n2000 = n961 | n1999 ;
  assign y0 = n85 ;
  assign y1 = n86 ;
  assign y2 = 1'b0 ;
  assign y3 = n87 ;
  assign y4 = n89 ;
  assign y5 = n116 ;
  assign y6 = n362 ;
  assign y7 = n367 ;
  assign y8 = n379 ;
  assign y9 = n381 ;
  assign y10 = n610 ;
  assign y11 = n681 ;
  assign y12 = n742 ;
  assign y13 = n840 ;
  assign y14 = n870 ;
  assign y15 = n1006 ;
  assign y16 = n1057 ;
  assign y17 = n1115 ;
  assign y18 = n1156 ;
  assign y19 = n1202 ;
  assign y20 = n428 ;
  assign y21 = n435 ;
  assign y22 = n1342 ;
  assign y23 = n1344 ;
  assign y24 = n1039 ;
  assign y25 = n1374 ;
  assign y26 = n1377 ;
  assign y27 = n1385 ;
  assign y28 = n1460 ;
  assign y29 = n1481 ;
  assign y30 = n1486 ;
  assign y31 = n1490 ;
  assign y32 = n1497 ;
  assign y33 = n1500 ;
  assign y34 = n1547 ;
  assign y35 = n1630 ;
  assign y36 = n1730 ;
  assign y37 = n1879 ;
  assign y38 = n1976 ;
  assign y39 = n1994 ;
  assign y40 = n2000 ;
  assign y41 = n264 ;
  assign y42 = 1'b0 ;
  assign y43 = n1331 ;
  assign y44 = n1039 ;
endmodule
