module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 ;
  assign n25 = x1 & x11 ;
  assign n26 = ( x0 & x10 ) | ( x0 & n25 ) | ( x10 & n25 ) ;
  assign n27 = ~x0 & n26 ;
  assign n28 = ( x1 & x9 ) | ( x1 & ~n27 ) | ( x9 & ~n27 ) ;
  assign n29 = x3 & n28 ;
  assign n30 = ( x3 & n27 ) | ( x3 & ~n29 ) | ( n27 & ~n29 ) ;
  assign n31 = ~x17 & x18 ;
  assign n32 = x16 & ~n31 ;
  assign n33 = ( x14 & ~n30 ) | ( x14 & n32 ) | ( ~n30 & n32 ) ;
  assign n34 = n30 & n33 ;
  assign n35 = ~x0 & x2 ;
  assign n36 = x1 & n35 ;
  assign n37 = x3 & n36 ;
  assign n38 = ( x5 & x18 ) | ( x5 & n37 ) | ( x18 & n37 ) ;
  assign n39 = ~x18 & n38 ;
  assign n40 = ( x2 & x5 ) | ( x2 & ~n39 ) | ( x5 & ~n39 ) ;
  assign n41 = n34 & n40 ;
  assign n42 = ( n34 & n39 ) | ( n34 & ~n41 ) | ( n39 & ~n41 ) ;
  assign n43 = ~x15 & n42 ;
  assign n44 = x1 & x3 ;
  assign n45 = ( x0 & x2 ) | ( x0 & n44 ) | ( x2 & n44 ) ;
  assign n46 = ~x0 & n45 ;
  assign n47 = x17 | x18 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = ( x5 & x15 ) | ( x5 & n48 ) | ( x15 & n48 ) ;
  assign n50 = ~x15 & n49 ;
  assign n51 = x14 & x16 ;
  assign n52 = x5 | x18 ;
  assign n53 = x9 | n52 ;
  assign n54 = ~x2 & x3 ;
  assign n55 = ( x1 & ~n53 ) | ( x1 & n54 ) | ( ~n53 & n54 ) ;
  assign n56 = ~x1 & n55 ;
  assign n57 = x10 & ~x18 ;
  assign n58 = x11 & n57 ;
  assign n59 = x3 & x17 ;
  assign n60 = ( ~x2 & x5 ) | ( ~x2 & n59 ) | ( x5 & n59 ) ;
  assign n61 = x2 & n60 ;
  assign n62 = ( x2 & x5 ) | ( x2 & ~n61 ) | ( x5 & ~n61 ) ;
  assign n63 = n58 & n62 ;
  assign n64 = ( n58 & n61 ) | ( n58 & ~n63 ) | ( n61 & ~n63 ) ;
  assign n65 = ( ~x0 & n56 ) | ( ~x0 & n64 ) | ( n56 & n64 ) ;
  assign n66 = x1 & ~n65 ;
  assign n67 = ( x1 & n56 ) | ( x1 & ~n66 ) | ( n56 & ~n66 ) ;
  assign n68 = ~x15 & n67 ;
  assign n69 = ( ~n51 & n67 ) | ( ~n51 & n68 ) | ( n67 & n68 ) ;
  assign n70 = n50 | n69 ;
  assign n71 = ( n42 & ~n43 ) | ( n42 & n70 ) | ( ~n43 & n70 ) ;
  assign n72 = x4 & n71 ;
  assign n73 = x1 & x5 ;
  assign n74 = ( x2 & n31 ) | ( x2 & n73 ) | ( n31 & n73 ) ;
  assign n75 = ~n31 & n74 ;
  assign n76 = ( x0 & x7 ) | ( x0 & n75 ) | ( x7 & n75 ) ;
  assign n77 = x1 | x9 ;
  assign n78 = x2 | n77 ;
  assign n79 = x7 & ~n78 ;
  assign n80 = ( ~x0 & n76 ) | ( ~x0 & n79 ) | ( n76 & n79 ) ;
  assign n81 = n72 | n80 ;
  assign n82 = ( x3 & n72 ) | ( x3 & n81 ) | ( n72 & n81 ) ;
  assign n83 = x13 & ~n82 ;
  assign n84 = ~x20 & x22 ;
  assign n85 = x21 & n84 ;
  assign n86 = ~x19 & n85 ;
  assign n87 = x13 | n86 ;
  assign n88 = ~n83 & n87 ;
  assign n89 = ~x3 & x14 ;
  assign n90 = x14 & ~x18 ;
  assign n91 = x3 & n90 ;
  assign n92 = ( x3 & n89 ) | ( x3 & ~n91 ) | ( n89 & ~n91 ) ;
  assign n93 = x16 & ~n92 ;
  assign n94 = x15 & n93 ;
  assign n95 = x15 & x16 ;
  assign n96 = ( x14 & x16 ) | ( x14 & n95 ) | ( x16 & n95 ) ;
  assign n97 = x14 & x15 ;
  assign n98 = ~x3 & n96 ;
  assign n99 = ( n96 & n97 ) | ( n96 & n98 ) | ( n97 & n98 ) ;
  assign n100 = ( x17 & ~n94 ) | ( x17 & n99 ) | ( ~n94 & n99 ) ;
  assign n101 = ~x18 & n100 ;
  assign n102 = ( x18 & ~n94 ) | ( x18 & n101 ) | ( ~n94 & n101 ) ;
  assign n103 = ( x4 & x5 ) | ( x4 & n102 ) | ( x5 & n102 ) ;
  assign n104 = x3 & ~x7 ;
  assign n105 = ~x3 & x6 ;
  assign n106 = ( x3 & ~n104 ) | ( x3 & n105 ) | ( ~n104 & n105 ) ;
  assign n107 = ( x17 & ~x18 ) | ( x17 & n106 ) | ( ~x18 & n106 ) ;
  assign n108 = ( x15 & ~x17 ) | ( x15 & n106 ) | ( ~x17 & n106 ) ;
  assign n109 = n107 & n108 ;
  assign n110 = x5 & n109 ;
  assign n111 = ( ~n102 & n103 ) | ( ~n102 & n110 ) | ( n103 & n110 ) ;
  assign n112 = x2 & ~n111 ;
  assign n113 = ( x16 & x17 ) | ( x16 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n114 = x14 & ~n113 ;
  assign n115 = ( ~x14 & x18 ) | ( ~x14 & n114 ) | ( x18 & n114 ) ;
  assign n116 = ( ~x11 & x15 ) | ( ~x11 & n115 ) | ( x15 & n115 ) ;
  assign n117 = ( x11 & x15 ) | ( x11 & ~x18 ) | ( x15 & ~x18 ) ;
  assign n118 = ~n116 & n117 ;
  assign n119 = x4 & x10 ;
  assign n120 = ( x5 & n118 ) | ( x5 & n119 ) | ( n118 & n119 ) ;
  assign n121 = ~x5 & n120 ;
  assign n122 = ~x2 & n121 ;
  assign n123 = ( x2 & ~n112 ) | ( x2 & n122 ) | ( ~n112 & n122 ) ;
  assign n124 = x1 & ~n123 ;
  assign n125 = ( x15 & x16 ) | ( x15 & ~n31 ) | ( x16 & ~n31 ) ;
  assign n126 = ( n31 & n51 ) | ( n31 & n125 ) | ( n51 & n125 ) ;
  assign n127 = ~x5 & x10 ;
  assign n128 = ( x4 & n126 ) | ( x4 & n127 ) | ( n126 & n127 ) ;
  assign n129 = ~n126 & n128 ;
  assign n130 = x2 & n129 ;
  assign n131 = x1 | n130 ;
  assign n132 = ~n124 & n131 ;
  assign n133 = ~x0 & n132 ;
  assign n134 = x3 & ~x9 ;
  assign n135 = ( ~x18 & n51 ) | ( ~x18 & n134 ) | ( n51 & n134 ) ;
  assign n136 = ~n51 & n135 ;
  assign n137 = x14 & ~n89 ;
  assign n138 = ~x9 & n137 ;
  assign n139 = ( x0 & ~n89 ) | ( x0 & n137 ) | ( ~n89 & n137 ) ;
  assign n140 = ( ~x3 & n138 ) | ( ~x3 & n139 ) | ( n138 & n139 ) ;
  assign n141 = ( ~n31 & n136 ) | ( ~n31 & n140 ) | ( n136 & n140 ) ;
  assign n142 = x16 & ~n141 ;
  assign n143 = ( x16 & n136 ) | ( x16 & ~n142 ) | ( n136 & ~n142 ) ;
  assign n144 = ( x5 & ~x15 ) | ( x5 & n143 ) | ( ~x15 & n143 ) ;
  assign n145 = x0 & ~n96 ;
  assign n146 = ~x3 & n145 ;
  assign n147 = x3 & ~x15 ;
  assign n148 = ( x9 & ~x18 ) | ( x9 & n147 ) | ( ~x18 & n147 ) ;
  assign n149 = ~x9 & n148 ;
  assign n150 = n146 | n149 ;
  assign n151 = ~x5 & n150 ;
  assign n152 = ( n143 & ~n144 ) | ( n143 & n151 ) | ( ~n144 & n151 ) ;
  assign n153 = ( x2 & ~x4 ) | ( x2 & n152 ) | ( ~x4 & n152 ) ;
  assign n154 = ~x6 & x9 ;
  assign n155 = x0 & ~x3 ;
  assign n156 = ( x6 & n154 ) | ( x6 & n155 ) | ( n154 & n155 ) ;
  assign n157 = x7 & n134 ;
  assign n158 = n156 | n157 ;
  assign n159 = ~x2 & n158 ;
  assign n160 = ( n152 & ~n153 ) | ( n152 & n159 ) | ( ~n153 & n159 ) ;
  assign n161 = n133 | n160 ;
  assign n162 = ( ~x1 & n133 ) | ( ~x1 & n161 ) | ( n133 & n161 ) ;
  assign n163 = x13 & n162 ;
  assign n164 = ( ~x19 & x20 ) | ( ~x19 & x22 ) | ( x20 & x22 ) ;
  assign n165 = ( ~x19 & x20 ) | ( ~x19 & x21 ) | ( x20 & x21 ) ;
  assign n166 = n164 & ~n165 ;
  assign n167 = x13 | n166 ;
  assign n168 = ( ~x13 & n163 ) | ( ~x13 & n167 ) | ( n163 & n167 ) ;
  assign n169 = ~x20 & n165 ;
  assign n170 = ( x21 & x22 ) | ( x21 & ~n169 ) | ( x22 & ~n169 ) ;
  assign n171 = ( n165 & n169 ) | ( n165 & ~n170 ) | ( n169 & ~n170 ) ;
  assign n172 = ~x13 & n171 ;
  assign n173 = x15 | x18 ;
  assign n174 = ( x18 & n51 ) | ( x18 & n173 ) | ( n51 & n173 ) ;
  assign n175 = ( x3 & ~x9 ) | ( x3 & n146 ) | ( ~x9 & n146 ) ;
  assign n176 = n174 | n175 ;
  assign n177 = ( n146 & ~n174 ) | ( n146 & n176 ) | ( ~n174 & n176 ) ;
  assign n178 = x4 & n177 ;
  assign n179 = ~x5 & n178 ;
  assign n180 = n158 & ~n179 ;
  assign n181 = x1 | x2 ;
  assign n182 = ( n179 & n180 ) | ( n179 & ~n181 ) | ( n180 & ~n181 ) ;
  assign n183 = ( ~x3 & x14 ) | ( ~x3 & x15 ) | ( x14 & x15 ) ;
  assign n184 = x16 & n183 ;
  assign n185 = ( x5 & x17 ) | ( x5 & n184 ) | ( x17 & n184 ) ;
  assign n186 = x3 & ~x17 ;
  assign n187 = ( ~x18 & n97 ) | ( ~x18 & n186 ) | ( n97 & n186 ) ;
  assign n188 = ~n97 & n187 ;
  assign n189 = x5 & n188 ;
  assign n190 = ( ~n184 & n185 ) | ( ~n184 & n189 ) | ( n185 & n189 ) ;
  assign n191 = x1 & n190 ;
  assign n192 = ~x1 & x5 ;
  assign n193 = x5 & ~n192 ;
  assign n194 = ~n47 & n193 ;
  assign n195 = ( x10 & ~n192 ) | ( x10 & n193 ) | ( ~n192 & n193 ) ;
  assign n196 = ( ~x1 & n194 ) | ( ~x1 & n195 ) | ( n194 & n195 ) ;
  assign n197 = n191 | n196 ;
  assign n198 = ( ~n96 & n191 ) | ( ~n96 & n197 ) | ( n191 & n197 ) ;
  assign n199 = x4 & n198 ;
  assign n200 = ~x15 & x17 ;
  assign n201 = ( x17 & n31 ) | ( x17 & ~n200 ) | ( n31 & ~n200 ) ;
  assign n202 = x5 & n106 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = n199 | n203 ;
  assign n205 = ( x1 & n199 ) | ( x1 & n204 ) | ( n199 & n204 ) ;
  assign n206 = ( x0 & ~x2 ) | ( x0 & n205 ) | ( ~x2 & n205 ) ;
  assign n207 = x11 & ~n174 ;
  assign n208 = ( x5 & x10 ) | ( x5 & n207 ) | ( x10 & n207 ) ;
  assign n209 = ~x5 & n208 ;
  assign n210 = x1 & x4 ;
  assign n211 = ( x2 & n209 ) | ( x2 & n210 ) | ( n209 & n210 ) ;
  assign n212 = ~x2 & n211 ;
  assign n213 = ~x0 & n212 ;
  assign n214 = ( n205 & ~n206 ) | ( n205 & n213 ) | ( ~n206 & n213 ) ;
  assign n215 = n182 | n214 ;
  assign n216 = x13 & n215 ;
  assign n217 = n172 | n216 ;
  assign n218 = ( x20 & x21 ) | ( x20 & x22 ) | ( x21 & x22 ) ;
  assign n219 = ~n164 & n218 ;
  assign n220 = x13 | n219 ;
  assign n221 = x3 & x11 ;
  assign n222 = x8 & n221 ;
  assign n223 = x0 & x1 ;
  assign n224 = x0 & ~n223 ;
  assign n225 = n222 & n224 ;
  assign n226 = ( x5 & n31 ) | ( x5 & n106 ) | ( n31 & n106 ) ;
  assign n227 = x3 | x14 ;
  assign n228 = x15 | n31 ;
  assign n229 = ( ~x3 & n227 ) | ( ~x3 & n228 ) | ( n227 & n228 ) ;
  assign n230 = ( ~x3 & x14 ) | ( ~x3 & n229 ) | ( x14 & n229 ) ;
  assign n231 = ~n47 & n230 ;
  assign n232 = ( n47 & n229 ) | ( n47 & n231 ) | ( n229 & n231 ) ;
  assign n233 = x16 | n201 ;
  assign n234 = ( x4 & n94 ) | ( x4 & ~n233 ) | ( n94 & ~n233 ) ;
  assign n235 = n232 & n234 ;
  assign n236 = ( x4 & ~n232 ) | ( x4 & n235 ) | ( ~n232 & n235 ) ;
  assign n237 = x5 & n236 ;
  assign n238 = ( ~n31 & n226 ) | ( ~n31 & n237 ) | ( n226 & n237 ) ;
  assign n239 = ( ~n223 & n224 ) | ( ~n223 & n238 ) | ( n224 & n238 ) ;
  assign n240 = ( x1 & n225 ) | ( x1 & n239 ) | ( n225 & n239 ) ;
  assign n241 = x2 & n240 ;
  assign n242 = x13 & ~n241 ;
  assign n243 = n220 & ~n242 ;
  assign n244 = ( x15 & x16 ) | ( x15 & x17 ) | ( x16 & x17 ) ;
  assign n245 = ( ~x17 & n51 ) | ( ~x17 & n244 ) | ( n51 & n244 ) ;
  assign n246 = ~x1 & x10 ;
  assign n247 = ( x2 & n245 ) | ( x2 & n246 ) | ( n245 & n246 ) ;
  assign n248 = ~n245 & n247 ;
  assign n249 = ( x0 & x13 ) | ( x0 & n248 ) | ( x13 & n248 ) ;
  assign n250 = ( x15 & ~x18 ) | ( x15 & n30 ) | ( ~x18 & n30 ) ;
  assign n251 = ~x14 & x16 ;
  assign n252 = ( x16 & x18 ) | ( x16 & ~n251 ) | ( x18 & ~n251 ) ;
  assign n253 = ( ~x16 & x17 ) | ( ~x16 & n251 ) | ( x17 & n251 ) ;
  assign n254 = ( ~x17 & n252 ) | ( ~x17 & n253 ) | ( n252 & n253 ) ;
  assign n255 = ( x15 & ~n30 ) | ( x15 & n254 ) | ( ~n30 & n254 ) ;
  assign n256 = n250 & ~n255 ;
  assign n257 = x0 & ~x1 ;
  assign n258 = ( ~x3 & n245 ) | ( ~x3 & n257 ) | ( n245 & n257 ) ;
  assign n259 = ~n245 & n258 ;
  assign n260 = ~x2 & n259 ;
  assign n261 = ( ~x2 & n256 ) | ( ~x2 & n260 ) | ( n256 & n260 ) ;
  assign n262 = x13 & n261 ;
  assign n263 = ( ~x0 & n249 ) | ( ~x0 & n262 ) | ( n249 & n262 ) ;
  assign n264 = x12 & x18 ;
  assign n265 = ( x4 & ~x5 ) | ( x4 & n264 ) | ( ~x5 & n264 ) ;
  assign n266 = n263 & ~n265 ;
  assign n267 = ( n263 & n264 ) | ( n263 & ~n266 ) | ( n264 & ~n266 ) ;
  assign n268 = x16 | x18 ;
  assign n269 = ( x16 & ~x17 ) | ( x16 & n268 ) | ( ~x17 & n268 ) ;
  assign n270 = ( x3 & ~n251 ) | ( x3 & n269 ) | ( ~n251 & n269 ) ;
  assign n271 = ( x14 & x18 ) | ( x14 & n31 ) | ( x18 & n31 ) ;
  assign n272 = ( ~x3 & n269 ) | ( ~x3 & n271 ) | ( n269 & n271 ) ;
  assign n273 = n270 & n272 ;
  assign n274 = ( x2 & n73 ) | ( x2 & n273 ) | ( n73 & n273 ) ;
  assign n275 = ~n273 & n274 ;
  assign n276 = ( x0 & x15 ) | ( x0 & n275 ) | ( x15 & n275 ) ;
  assign n277 = ~x2 & n140 ;
  assign n278 = ~x1 & n277 ;
  assign n279 = ~x1 & x2 ;
  assign n280 = x1 & x14 ;
  assign n281 = ~x2 & x11 ;
  assign n282 = x14 & ~n281 ;
  assign n283 = ( n279 & n280 ) | ( n279 & ~n282 ) | ( n280 & ~n282 ) ;
  assign n284 = ( ~x0 & n278 ) | ( ~x0 & n283 ) | ( n278 & n283 ) ;
  assign n285 = x10 & ~n284 ;
  assign n286 = ( x10 & n278 ) | ( x10 & ~n285 ) | ( n278 & ~n285 ) ;
  assign n287 = ~n31 & n286 ;
  assign n288 = ( x5 & ~x16 ) | ( x5 & n287 ) | ( ~x16 & n287 ) ;
  assign n289 = ( x1 & ~x16 ) | ( x1 & n155 ) | ( ~x16 & n155 ) ;
  assign n290 = ~x1 & n289 ;
  assign n291 = ~x18 & n30 ;
  assign n292 = ~n51 & n291 ;
  assign n293 = x2 & ~x16 ;
  assign n294 = x10 & n293 ;
  assign n295 = ~x0 & n294 ;
  assign n296 = ~x1 & n295 ;
  assign n297 = ( ~n290 & n292 ) | ( ~n290 & n296 ) | ( n292 & n296 ) ;
  assign n298 = x2 & ~n296 ;
  assign n299 = ( n290 & n297 ) | ( n290 & ~n298 ) | ( n297 & ~n298 ) ;
  assign n300 = ~x5 & n299 ;
  assign n301 = ( n287 & ~n288 ) | ( n287 & n300 ) | ( ~n288 & n300 ) ;
  assign n302 = x15 & n301 ;
  assign n303 = ( ~x0 & n276 ) | ( ~x0 & n302 ) | ( n276 & n302 ) ;
  assign n304 = ( x4 & n264 ) | ( x4 & n303 ) | ( n264 & n303 ) ;
  assign n305 = x13 & ~n304 ;
  assign n306 = ( x13 & n264 ) | ( x13 & ~n305 ) | ( n264 & ~n305 ) ;
  assign n307 = ( ~x3 & x6 ) | ( ~x3 & x8 ) | ( x6 & x8 ) ;
  assign n308 = ~x9 & n307 ;
  assign n309 = ( ~x3 & x9 ) | ( ~x3 & n308 ) | ( x9 & n308 ) ;
  assign n310 = x0 | n157 ;
  assign n311 = ( n157 & n309 ) | ( n157 & n310 ) | ( n309 & n310 ) ;
  assign n312 = ~x1 & x13 ;
  assign n313 = ( x2 & n311 ) | ( x2 & ~n312 ) | ( n311 & ~n312 ) ;
  assign n314 = n311 & ~n313 ;
  assign n315 = ( x16 & n47 ) | ( x16 & n51 ) | ( n47 & n51 ) ;
  assign n316 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n317 = x14 & ~n316 ;
  assign n318 = ( x14 & x18 ) | ( x14 & ~n317 ) | ( x18 & ~n317 ) ;
  assign n319 = x9 | n318 ;
  assign n320 = ( x2 & x3 ) | ( x2 & ~n319 ) | ( x3 & ~n319 ) ;
  assign n321 = ~x2 & n320 ;
  assign n322 = x0 & x2 ;
  assign n323 = x2 & ~n322 ;
  assign n324 = x10 & n323 ;
  assign n325 = ( x3 & n322 ) | ( x3 & ~n323 ) | ( n322 & ~n323 ) ;
  assign n326 = ( x0 & n324 ) | ( x0 & ~n325 ) | ( n324 & ~n325 ) ;
  assign n327 = n321 | n326 ;
  assign n328 = ( ~n315 & n321 ) | ( ~n315 & n327 ) | ( n321 & n327 ) ;
  assign n329 = x1 | n328 ;
  assign n330 = x11 & ~n318 ;
  assign n331 = ( x2 & x10 ) | ( x2 & n330 ) | ( x10 & n330 ) ;
  assign n332 = ~x2 & n331 ;
  assign n333 = ~x0 & n332 ;
  assign n334 = x1 & ~n333 ;
  assign n335 = n329 & ~n334 ;
  assign n336 = ~x5 & x15 ;
  assign n337 = ( x13 & ~n335 ) | ( x13 & n336 ) | ( ~n335 & n336 ) ;
  assign n338 = n335 & n337 ;
  assign n339 = n264 | n338 ;
  assign n340 = ( x4 & n264 ) | ( x4 & n339 ) | ( n264 & n339 ) ;
  assign n341 = ( x5 & ~x6 ) | ( x5 & n96 ) | ( ~x6 & n96 ) ;
  assign n342 = x4 & n341 ;
  assign n343 = ( x4 & x6 ) | ( x4 & ~n342 ) | ( x6 & ~n342 ) ;
  assign n344 = ( x1 & ~x2 ) | ( x1 & n343 ) | ( ~x2 & n343 ) ;
  assign n345 = ~x2 & x8 ;
  assign n346 = ( ~x1 & n344 ) | ( ~x1 & n345 ) | ( n344 & n345 ) ;
  assign n347 = x0 & n346 ;
  assign n348 = x6 & ~n47 ;
  assign n349 = x5 & n348 ;
  assign n350 = n347 | n349 ;
  assign n351 = ( n36 & n347 ) | ( n36 & n350 ) | ( n347 & n350 ) ;
  assign n352 = ( x3 & ~x13 ) | ( x3 & n351 ) | ( ~x13 & n351 ) ;
  assign n353 = x5 & ~n47 ;
  assign n354 = n36 & n353 ;
  assign n355 = ~x15 & n51 ;
  assign n356 = x5 | x9 ;
  assign n357 = ( n51 & ~n355 ) | ( n51 & n356 ) | ( ~n355 & n356 ) ;
  assign n358 = x5 & ~n97 ;
  assign n359 = ~x17 & n358 ;
  assign n360 = x2 & n359 ;
  assign n361 = ( x0 & x1 ) | ( x0 & n360 ) | ( x1 & n360 ) ;
  assign n362 = ~x0 & n361 ;
  assign n363 = ( x1 & x2 ) | ( x1 & ~n362 ) | ( x2 & ~n362 ) ;
  assign n364 = ~n357 & n363 ;
  assign n365 = ( n357 & ~n362 ) | ( n357 & n364 ) | ( ~n362 & n364 ) ;
  assign n366 = ( x4 & ~x18 ) | ( x4 & n365 ) | ( ~x18 & n365 ) ;
  assign n367 = x23 & ~n97 ;
  assign n368 = x5 & n367 ;
  assign n369 = x2 & n368 ;
  assign n370 = ( x0 & x1 ) | ( x0 & n369 ) | ( x1 & n369 ) ;
  assign n371 = ~x0 & n370 ;
  assign n372 = ~x18 & n371 ;
  assign n373 = ( ~n365 & n366 ) | ( ~n365 & n372 ) | ( n366 & n372 ) ;
  assign n374 = ( n78 & n354 ) | ( n78 & ~n373 ) | ( n354 & ~n373 ) ;
  assign n375 = x7 | n373 ;
  assign n376 = ( n354 & ~n374 ) | ( n354 & n375 ) | ( ~n374 & n375 ) ;
  assign n377 = x3 & n376 ;
  assign n378 = ( x1 & x4 ) | ( x1 & n127 ) | ( x4 & n127 ) ;
  assign n379 = ~x1 & n378 ;
  assign n380 = ( x4 & x17 ) | ( x4 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n381 = ~x18 & x23 ;
  assign n382 = ( ~x17 & n380 ) | ( ~x17 & n381 ) | ( n380 & n381 ) ;
  assign n383 = ( x1 & n379 ) | ( x1 & n382 ) | ( n379 & n382 ) ;
  assign n384 = x5 & ~n383 ;
  assign n385 = ( x5 & n379 ) | ( x5 & ~n384 ) | ( n379 & ~n384 ) ;
  assign n386 = ( ~n96 & n212 ) | ( ~n96 & n385 ) | ( n212 & n385 ) ;
  assign n387 = x2 & ~n386 ;
  assign n388 = ( x2 & n212 ) | ( x2 & ~n387 ) | ( n212 & ~n387 ) ;
  assign n389 = n377 | n388 ;
  assign n390 = ( ~x0 & n377 ) | ( ~x0 & n389 ) | ( n377 & n389 ) ;
  assign n391 = x13 & n390 ;
  assign n392 = ( n351 & ~n352 ) | ( n351 & n391 ) | ( ~n352 & n391 ) ;
  assign n393 = ( x3 & x14 ) | ( x3 & x17 ) | ( x14 & x17 ) ;
  assign n394 = ~x16 & x17 ;
  assign n395 = ( ~x14 & n393 ) | ( ~x14 & n394 ) | ( n393 & n394 ) ;
  assign n396 = ( x2 & n73 ) | ( x2 & ~n395 ) | ( n73 & ~n395 ) ;
  assign n397 = n395 & n396 ;
  assign n398 = ( x0 & x4 ) | ( x0 & n397 ) | ( x4 & n397 ) ;
  assign n399 = ( x5 & x16 ) | ( x5 & n287 ) | ( x16 & n287 ) ;
  assign n400 = x5 & ~n92 ;
  assign n401 = x2 & n400 ;
  assign n402 = ( x0 & x1 ) | ( x0 & n401 ) | ( x1 & n401 ) ;
  assign n403 = ~x0 & n402 ;
  assign n404 = x16 & n403 ;
  assign n405 = ( ~x5 & n399 ) | ( ~x5 & n404 ) | ( n399 & n404 ) ;
  assign n406 = x4 & n405 ;
  assign n407 = ( ~x0 & n398 ) | ( ~x0 & n406 ) | ( n398 & n406 ) ;
  assign n408 = ( x3 & ~x7 ) | ( x3 & x17 ) | ( ~x7 & x17 ) ;
  assign n409 = n51 & n381 ;
  assign n410 = x3 & n409 ;
  assign n411 = ( x7 & n408 ) | ( x7 & n410 ) | ( n408 & n410 ) ;
  assign n412 = ( x3 & x6 ) | ( x3 & ~x17 ) | ( x6 & ~x17 ) ;
  assign n413 = n251 & n381 ;
  assign n414 = ~x3 & n413 ;
  assign n415 = ( x6 & ~n412 ) | ( x6 & n414 ) | ( ~n412 & n414 ) ;
  assign n416 = ~n411 & n415 ;
  assign n417 = x2 & x5 ;
  assign n418 = ( n411 & n416 ) | ( n411 & n417 ) | ( n416 & n417 ) ;
  assign n419 = ( ~x0 & n407 ) | ( ~x0 & n418 ) | ( n407 & n418 ) ;
  assign n420 = x1 & ~n419 ;
  assign n421 = ( x1 & n407 ) | ( x1 & ~n420 ) | ( n407 & ~n420 ) ;
  assign n422 = ( x13 & x15 ) | ( x13 & ~n421 ) | ( x15 & ~n421 ) ;
  assign n423 = x4 & ~n51 ;
  assign n424 = x6 | n423 ;
  assign n425 = ( ~x3 & n423 ) | ( ~x3 & n424 ) | ( n423 & n424 ) ;
  assign n426 = ( ~x4 & x7 ) | ( ~x4 & n425 ) | ( x7 & n425 ) ;
  assign n427 = x3 | n425 ;
  assign n428 = ( x4 & n426 ) | ( x4 & n427 ) | ( n426 & n427 ) ;
  assign n429 = ( x5 & n200 ) | ( x5 & ~n428 ) | ( n200 & ~n428 ) ;
  assign n430 = n428 & n429 ;
  assign n431 = x2 & n430 ;
  assign n432 = ( x0 & x1 ) | ( x0 & n431 ) | ( x1 & n431 ) ;
  assign n433 = ~x0 & n432 ;
  assign n434 = x13 & n433 ;
  assign n435 = ( n421 & n422 ) | ( n421 & n434 ) | ( n422 & n434 ) ;
  assign n436 = ( ~x18 & n51 ) | ( ~x18 & n281 ) | ( n51 & n281 ) ;
  assign n437 = ~n51 & n436 ;
  assign n438 = ( x1 & x15 ) | ( x1 & ~n437 ) | ( x15 & ~n437 ) ;
  assign n439 = n32 & n283 ;
  assign n440 = x15 & n439 ;
  assign n441 = ( n437 & n438 ) | ( n437 & n440 ) | ( n438 & n440 ) ;
  assign n442 = x11 & ~x15 ;
  assign n443 = ~x18 & n442 ;
  assign n444 = x1 & x2 ;
  assign n445 = x1 & ~n444 ;
  assign n446 = n443 & n445 ;
  assign n447 = ( n96 & n444 ) | ( n96 & ~n445 ) | ( n444 & ~n445 ) ;
  assign n448 = ( x2 & n446 ) | ( x2 & ~n447 ) | ( n446 & ~n447 ) ;
  assign n449 = ~n441 & n448 ;
  assign n450 = x10 & x13 ;
  assign n451 = ( n441 & n449 ) | ( n441 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ~x5 & n451 ;
  assign n453 = ( x0 & x4 ) | ( x0 & n452 ) | ( x4 & n452 ) ;
  assign n454 = ~x0 & n453 ;
  assign n455 = x0 & ~x2 ;
  assign n456 = ( x1 & ~x3 ) | ( x1 & n455 ) | ( ~x3 & n455 ) ;
  assign n457 = ~x1 & n456 ;
  assign n458 = x13 & n457 ;
  assign n459 = x9 & n458 ;
  assign n460 = ( x1 & x2 ) | ( x1 & ~x13 ) | ( x2 & ~x13 ) ;
  assign n461 = ( x2 & ~x3 ) | ( x2 & x13 ) | ( ~x3 & x13 ) ;
  assign n462 = ~n460 & n461 ;
  assign n463 = x8 & n462 ;
  assign n464 = x0 & n463 ;
  assign n465 = x15 & ~x17 ;
  assign n466 = ( x5 & ~x18 ) | ( x5 & n465 ) | ( ~x18 & n465 ) ;
  assign n467 = ~x5 & n466 ;
  assign y0 = n88 ;
  assign y1 = n168 ;
  assign y2 = n217 ;
  assign y3 = n243 ;
  assign y4 = n267 ;
  assign y5 = n306 ;
  assign y6 = n314 ;
  assign y7 = n340 ;
  assign y8 = n392 ;
  assign y9 = n435 ;
  assign y10 = n454 ;
  assign y11 = n459 ;
  assign y12 = n464 ;
  assign y13 = n467 ;
endmodule
