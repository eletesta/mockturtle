module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 ;
  assign n34 = ( x9 & ~x11 ) | ( x9 & x14 ) | ( ~x11 & x14 ) ;
  assign n35 = ( ~x9 & x11 ) | ( ~x9 & n34 ) | ( x11 & n34 ) ;
  assign n36 = ( ~x14 & n34 ) | ( ~x14 & n35 ) | ( n34 & n35 ) ;
  assign n37 = ( x2 & x5 ) | ( x2 & n36 ) | ( x5 & n36 ) ;
  assign n38 = ( x2 & n36 ) | ( x2 & ~n37 ) | ( n36 & ~n37 ) ;
  assign n39 = ( x5 & ~n37 ) | ( x5 & n38 ) | ( ~n37 & n38 ) ;
  assign n40 = ~x7 & n39 ;
  assign n41 = x7 & ~n39 ;
  assign n42 = n40 | n41 ;
  assign n43 = x18 & ~x32 ;
  assign n44 = x22 & n43 ;
  assign n45 = n42 | n44 ;
  assign n46 = n42 & n44 ;
  assign n47 = n45 & ~n46 ;
  assign n48 = x30 & n47 ;
  assign n49 = ( x27 & n47 ) | ( x27 & n48 ) | ( n47 & n48 ) ;
  assign n50 = ( x27 & ~n47 ) | ( x27 & n48 ) | ( ~n47 & n48 ) ;
  assign n51 = ( n47 & ~n49 ) | ( n47 & n50 ) | ( ~n49 & n50 ) ;
  assign n52 = ( x1 & ~x4 ) | ( x1 & x7 ) | ( ~x4 & x7 ) ;
  assign n53 = ( ~x1 & x4 ) | ( ~x1 & n52 ) | ( x4 & n52 ) ;
  assign n54 = ( ~x7 & n52 ) | ( ~x7 & n53 ) | ( n52 & n53 ) ;
  assign n55 = ( x8 & ~x13 ) | ( x8 & x15 ) | ( ~x13 & x15 ) ;
  assign n56 = ( ~x8 & x13 ) | ( ~x8 & n55 ) | ( x13 & n55 ) ;
  assign n57 = ( ~x15 & n55 ) | ( ~x15 & n56 ) | ( n55 & n56 ) ;
  assign n58 = x23 | x32 ;
  assign n59 = x17 & ~n58 ;
  assign n60 = x14 & ~n59 ;
  assign n61 = ~x14 & n59 ;
  assign n62 = n60 | n61 ;
  assign n63 = ( n54 & n57 ) | ( n54 & n62 ) | ( n57 & n62 ) ;
  assign n64 = ( n57 & n62 ) | ( n57 & ~n63 ) | ( n62 & ~n63 ) ;
  assign n65 = ( n54 & ~n63 ) | ( n54 & n64 ) | ( ~n63 & n64 ) ;
  assign n66 = ~x10 & n65 ;
  assign n67 = x10 & ~n65 ;
  assign n68 = n66 | n67 ;
  assign n69 = x30 & n68 ;
  assign n70 = ( x26 & n68 ) | ( x26 & n69 ) | ( n68 & n69 ) ;
  assign n71 = ( x26 & ~n68 ) | ( x26 & n69 ) | ( ~n68 & n69 ) ;
  assign n72 = ( n68 & ~n70 ) | ( n68 & n71 ) | ( ~n70 & n71 ) ;
  assign n73 = n51 | n72 ;
  assign n74 = x22 & ~x23 ;
  assign n75 = x31 & ~x32 ;
  assign n76 = ( ~x22 & n74 ) | ( ~x22 & n75 ) | ( n74 & n75 ) ;
  assign n77 = ~x23 & x32 ;
  assign n78 = ( ~x22 & x32 ) | ( ~x22 & n77 ) | ( x32 & n77 ) ;
  assign n79 = ( ~x28 & n76 ) | ( ~x28 & n78 ) | ( n76 & n78 ) ;
  assign n80 = x30 & ~n79 ;
  assign n81 = ( x30 & n76 ) | ( x30 & ~n80 ) | ( n76 & ~n80 ) ;
  assign n82 = x16 & x30 ;
  assign n83 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n84 = ( ~x0 & x1 ) | ( ~x0 & n83 ) | ( x1 & n83 ) ;
  assign n85 = ( ~x2 & n83 ) | ( ~x2 & n84 ) | ( n83 & n84 ) ;
  assign n86 = ( x4 & x5 ) | ( x4 & n85 ) | ( x5 & n85 ) ;
  assign n87 = ( x4 & n85 ) | ( x4 & ~n86 ) | ( n85 & ~n86 ) ;
  assign n88 = ( x5 & ~n86 ) | ( x5 & n87 ) | ( ~n86 & n87 ) ;
  assign n89 = ~x6 & n88 ;
  assign n90 = x6 & ~n88 ;
  assign n91 = n89 | n90 ;
  assign n92 = ( ~x3 & x7 ) | ( ~x3 & n91 ) | ( x7 & n91 ) ;
  assign n93 = ( x3 & ~n91 ) | ( x3 & n92 ) | ( ~n91 & n92 ) ;
  assign n94 = ( ~x7 & n92 ) | ( ~x7 & n93 ) | ( n92 & n93 ) ;
  assign n95 = ( x9 & ~x14 ) | ( x9 & x15 ) | ( ~x14 & x15 ) ;
  assign n96 = ( ~x9 & x14 ) | ( ~x9 & n95 ) | ( x14 & n95 ) ;
  assign n97 = ( ~x15 & n95 ) | ( ~x15 & n96 ) | ( n95 & n96 ) ;
  assign n98 = x20 & ~x32 ;
  assign n99 = ( x8 & n97 ) | ( x8 & ~n98 ) | ( n97 & ~n98 ) ;
  assign n100 = ( ~n97 & n98 ) | ( ~n97 & n99 ) | ( n98 & n99 ) ;
  assign n101 = ( ~x8 & n99 ) | ( ~x8 & n100 ) | ( n99 & n100 ) ;
  assign n102 = ~n94 & n101 ;
  assign n103 = n94 & n101 ;
  assign n104 = ( n94 & n102 ) | ( n94 & ~n103 ) | ( n102 & ~n103 ) ;
  assign n105 = ( x16 & x23 ) | ( x16 & x30 ) | ( x23 & x30 ) ;
  assign n106 = n104 & n105 ;
  assign n107 = ( ~x30 & n104 ) | ( ~x30 & n105 ) | ( n104 & n105 ) ;
  assign n108 = ( n82 & ~n106 ) | ( n82 & n107 ) | ( ~n106 & n107 ) ;
  assign n109 = x17 & x30 ;
  assign n110 = ( x17 & x23 ) | ( x17 & n109 ) | ( x23 & n109 ) ;
  assign n111 = x21 & ~x32 ;
  assign n112 = ( x3 & x13 ) | ( x3 & ~n111 ) | ( x13 & ~n111 ) ;
  assign n113 = ( ~x3 & n111 ) | ( ~x3 & n112 ) | ( n111 & n112 ) ;
  assign n114 = ( ~x13 & n112 ) | ( ~x13 & n113 ) | ( n112 & n113 ) ;
  assign n115 = ( x10 & ~x11 ) | ( x10 & x12 ) | ( ~x11 & x12 ) ;
  assign n116 = ( ~x10 & x11 ) | ( ~x10 & n115 ) | ( x11 & n115 ) ;
  assign n117 = ( ~x12 & n115 ) | ( ~x12 & n116 ) | ( n115 & n116 ) ;
  assign n118 = ( n85 & n97 ) | ( n85 & n117 ) | ( n97 & n117 ) ;
  assign n119 = ( n97 & n117 ) | ( n97 & ~n118 ) | ( n117 & ~n118 ) ;
  assign n120 = ( n85 & ~n118 ) | ( n85 & n119 ) | ( ~n118 & n119 ) ;
  assign n121 = n114 & n120 ;
  assign n122 = n114 | n120 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = x30 & n123 ;
  assign n125 = ( x24 & n123 ) | ( x24 & n124 ) | ( n123 & n124 ) ;
  assign n126 = ( x24 & ~n123 ) | ( x24 & n124 ) | ( ~n123 & n124 ) ;
  assign n127 = ( n123 & ~n125 ) | ( n123 & n126 ) | ( ~n125 & n126 ) ;
  assign n128 = x19 & x30 ;
  assign n129 = ( x19 & ~x22 ) | ( x19 & n128 ) | ( ~x22 & n128 ) ;
  assign n130 = n127 & ~n129 ;
  assign n131 = ( n108 & n110 ) | ( n108 & ~n130 ) | ( n110 & ~n130 ) ;
  assign n132 = n108 & ~n131 ;
  assign n133 = n97 & ~n117 ;
  assign n134 = n97 | n117 ;
  assign n135 = ( ~n97 & n133 ) | ( ~n97 & n134 ) | ( n133 & n134 ) ;
  assign n136 = ( x4 & x5 ) | ( x4 & n135 ) | ( x5 & n135 ) ;
  assign n137 = ( x4 & n135 ) | ( x4 & ~n136 ) | ( n135 & ~n136 ) ;
  assign n138 = ( x5 & ~n136 ) | ( x5 & n137 ) | ( ~n136 & n137 ) ;
  assign n139 = ~x6 & n138 ;
  assign n140 = x6 & ~n138 ;
  assign n141 = n139 | n140 ;
  assign n142 = x16 & ~n58 ;
  assign n143 = x0 & ~n142 ;
  assign n144 = ~x0 & n142 ;
  assign n145 = n143 | n144 ;
  assign n146 = ( x25 & n141 ) | ( x25 & n145 ) | ( n141 & n145 ) ;
  assign n147 = ~x30 & n146 ;
  assign n148 = ( n141 & n145 ) | ( n141 & ~n146 ) | ( n145 & ~n146 ) ;
  assign n149 = ~x30 & n148 ;
  assign n150 = ( x25 & ~n147 ) | ( x25 & n149 ) | ( ~n147 & n149 ) ;
  assign n151 = x18 & x30 ;
  assign n152 = ( x3 & x6 ) | ( x3 & n57 ) | ( x6 & n57 ) ;
  assign n153 = ( x3 & n57 ) | ( x3 & ~n152 ) | ( n57 & ~n152 ) ;
  assign n154 = ( x6 & ~n152 ) | ( x6 & n153 ) | ( ~n152 & n153 ) ;
  assign n155 = ~x9 & n154 ;
  assign n156 = x9 & ~n154 ;
  assign n157 = n155 | n156 ;
  assign n158 = x19 & ~x32 ;
  assign n159 = x22 & n158 ;
  assign n160 = x12 & ~n159 ;
  assign n161 = ~x12 & n159 ;
  assign n162 = n160 | n161 ;
  assign n163 = n157 | n162 ;
  assign n164 = n157 & ~n162 ;
  assign n165 = ( ~n157 & n163 ) | ( ~n157 & n164 ) | ( n163 & n164 ) ;
  assign n166 = ( x18 & ~x22 ) | ( x18 & x30 ) | ( ~x22 & x30 ) ;
  assign n167 = n165 & n166 ;
  assign n168 = ( ~x30 & n165 ) | ( ~x30 & n166 ) | ( n165 & n166 ) ;
  assign n169 = ( n151 & ~n167 ) | ( n151 & n168 ) | ( ~n167 & n168 ) ;
  assign n170 = n150 & ~n169 ;
  assign n171 = n132 & n170 ;
  assign n172 = n81 & n171 ;
  assign n173 = ~n73 & n172 ;
  assign n174 = x0 & ~n173 ;
  assign n175 = ~x0 & n173 ;
  assign n176 = n174 | n175 ;
  assign n177 = ~n51 & n72 ;
  assign n178 = n150 | n169 ;
  assign n179 = n132 & ~n178 ;
  assign n180 = n81 & n179 ;
  assign n181 = n177 & n180 ;
  assign n182 = x1 & ~n181 ;
  assign n183 = ~x1 & n181 ;
  assign n184 = n182 | n183 ;
  assign n185 = n51 & ~n72 ;
  assign n186 = n180 & n185 ;
  assign n187 = x2 & ~n186 ;
  assign n188 = ~x2 & n186 ;
  assign n189 = n187 | n188 ;
  assign n190 = ~n150 & n169 ;
  assign n191 = n132 & n190 ;
  assign n192 = n81 & n191 ;
  assign n193 = ~n73 & n192 ;
  assign n194 = x3 & ~n193 ;
  assign n195 = ~x3 & n193 ;
  assign n196 = n194 | n195 ;
  assign n197 = ( ~x29 & n76 ) | ( ~x29 & n78 ) | ( n76 & n78 ) ;
  assign n198 = x30 & ~n197 ;
  assign n199 = ( x30 & n76 ) | ( x30 & ~n198 ) | ( n76 & ~n198 ) ;
  assign n200 = n150 & n169 ;
  assign n201 = n132 & n200 ;
  assign n202 = n199 & n201 ;
  assign n203 = n185 & n202 ;
  assign n204 = x9 & ~n203 ;
  assign n205 = ~x9 & n203 ;
  assign n206 = n204 | n205 ;
  assign n207 = n51 & n72 ;
  assign n208 = n171 & n199 ;
  assign n209 = n207 & n208 ;
  assign n210 = x14 & ~n209 ;
  assign n211 = ~x14 & n209 ;
  assign n212 = n210 | n211 ;
  assign n213 = n177 & n202 ;
  assign n214 = x15 & ~n213 ;
  assign n215 = ~x15 & n213 ;
  assign n216 = n214 | n215 ;
  assign n217 = n127 | n129 ;
  assign n218 = n108 & ~n217 ;
  assign n219 = ~n110 & n218 ;
  assign n220 = n170 & n219 ;
  assign n221 = n81 & n220 ;
  assign n222 = n177 & n221 ;
  assign n223 = x4 & ~n222 ;
  assign n224 = ~x4 & n222 ;
  assign n225 = n223 | n224 ;
  assign n226 = n185 & n221 ;
  assign n227 = x5 & ~n226 ;
  assign n228 = ~x5 & n226 ;
  assign n229 = n227 | n228 ;
  assign n230 = n200 & n219 ;
  assign n231 = n81 & n230 ;
  assign n232 = ~n73 & n231 ;
  assign n233 = x6 & ~n232 ;
  assign n234 = ~x6 & n232 ;
  assign n235 = n233 | n234 ;
  assign n236 = ~n178 & n219 ;
  assign n237 = n81 & n236 ;
  assign n238 = n207 & n237 ;
  assign n239 = x7 & ~n238 ;
  assign n240 = ~x7 & n238 ;
  assign n241 = n239 | n240 ;
  assign n242 = n190 & n219 ;
  assign n243 = n199 & n242 ;
  assign n244 = n177 & n243 ;
  assign n245 = x8 & ~n244 ;
  assign n246 = ~x8 & n244 ;
  assign n247 = n245 | n246 ;
  assign n248 = n108 | n110 ;
  assign n249 = n127 & ~n248 ;
  assign n250 = ~n129 & n249 ;
  assign n251 = n170 & n250 ;
  assign n252 = n199 & n251 ;
  assign n253 = n177 & n252 ;
  assign n254 = x10 & ~n253 ;
  assign n255 = ~x10 & n253 ;
  assign n256 = n254 | n255 ;
  assign n257 = n185 & n252 ;
  assign n258 = x11 & ~n257 ;
  assign n259 = ~x11 & n257 ;
  assign n260 = n258 | n259 ;
  assign n261 = n200 & n250 ;
  assign n262 = n199 & n261 ;
  assign n263 = ~n73 & n262 ;
  assign n264 = x12 & ~n263 ;
  assign n265 = ~x12 & n263 ;
  assign n266 = n264 | n265 ;
  assign n267 = n177 & n250 ;
  assign n268 = ( n190 & ~n199 ) | ( n190 & n267 ) | ( ~n199 & n267 ) ;
  assign n269 = n199 & n268 ;
  assign n270 = ~x13 & n269 ;
  assign n271 = x13 | n269 ;
  assign n272 = ( ~n269 & n270 ) | ( ~n269 & n271 ) | ( n270 & n271 ) ;
  assign n273 = n217 | n248 ;
  assign n274 = n190 & ~n273 ;
  assign n275 = n129 & ~n178 ;
  assign n276 = ( ~n127 & n248 ) | ( ~n127 & n275 ) | ( n248 & n275 ) ;
  assign n277 = ~n248 & n276 ;
  assign n278 = n76 & n177 ;
  assign n279 = ( ~n178 & n273 ) | ( ~n178 & n278 ) | ( n273 & n278 ) ;
  assign n280 = ~n273 & n279 ;
  assign n281 = n76 & ~n178 ;
  assign n282 = ( n185 & n273 ) | ( n185 & n281 ) | ( n273 & n281 ) ;
  assign n283 = ~n273 & n282 ;
  assign n284 = n219 & ~n250 ;
  assign n285 = ~n73 & n76 ;
  assign n286 = ~n178 & n285 ;
  assign n287 = ( n250 & n284 ) | ( n250 & n286 ) | ( n284 & n286 ) ;
  assign n288 = ( ~n273 & n285 ) | ( ~n273 & n287 ) | ( n285 & n287 ) ;
  assign n289 = n170 & ~n288 ;
  assign n290 = ( n170 & n287 ) | ( n170 & ~n289 ) | ( n287 & ~n289 ) ;
  assign n291 = n283 | n290 ;
  assign n292 = n280 | n291 ;
  assign n293 = ( ~n274 & n277 ) | ( ~n274 & n292 ) | ( n277 & n292 ) ;
  assign n294 = n285 | n292 ;
  assign n295 = ( n274 & n293 ) | ( n274 & n294 ) | ( n293 & n294 ) ;
  assign n296 = ~n108 & n110 ;
  assign n297 = ~n217 & n296 ;
  assign n298 = ( n178 & n285 ) | ( n178 & ~n297 ) | ( n285 & ~n297 ) ;
  assign n299 = n285 & ~n298 ;
  assign n300 = n177 & n199 ;
  assign n301 = n201 & ~n300 ;
  assign n302 = ( ~n73 & n81 ) | ( ~n73 & n181 ) | ( n81 & n181 ) ;
  assign n303 = n171 & ~n302 ;
  assign n304 = ( n171 & n181 ) | ( n171 & ~n303 ) | ( n181 & ~n303 ) ;
  assign n305 = n193 | n304 ;
  assign n306 = ( n186 & ~n222 ) | ( n186 & n305 ) | ( ~n222 & n305 ) ;
  assign n307 = n222 | n306 ;
  assign n308 = n232 | n307 ;
  assign n309 = ( n226 & ~n238 ) | ( n226 & n308 ) | ( ~n238 & n308 ) ;
  assign n310 = n238 | n309 ;
  assign n311 = n190 & n250 ;
  assign n312 = n300 & n311 ;
  assign n313 = n185 & n199 ;
  assign n314 = n201 & n313 ;
  assign n315 = n242 | n314 ;
  assign n316 = ( n300 & n314 ) | ( n300 & n315 ) | ( n314 & n315 ) ;
  assign n317 = ( ~n300 & n313 ) | ( ~n300 & n316 ) | ( n313 & n316 ) ;
  assign n318 = n251 | n316 ;
  assign n319 = ( n300 & n317 ) | ( n300 & n318 ) | ( n317 & n318 ) ;
  assign n320 = n209 | n319 ;
  assign n321 = ( ~n263 & n312 ) | ( ~n263 & n320 ) | ( n312 & n320 ) ;
  assign n322 = n263 | n321 ;
  assign n323 = n310 | n322 ;
  assign n324 = ( n201 & ~n301 ) | ( n201 & n323 ) | ( ~n301 & n323 ) ;
  assign n325 = n299 | n324 ;
  assign n326 = n295 | n325 ;
  assign n327 = ~x31 & n326 ;
  assign n328 = n110 | n127 ;
  assign n329 = n72 | n169 ;
  assign n330 = ( ~n51 & n150 ) | ( ~n51 & n329 ) | ( n150 & n329 ) ;
  assign n331 = n51 | n330 ;
  assign n332 = n108 | n331 ;
  assign n333 = ( ~n129 & n328 ) | ( ~n129 & n332 ) | ( n328 & n332 ) ;
  assign n334 = n129 | n333 ;
  assign n335 = ~x32 & n334 ;
  assign n336 = ( ~n326 & n327 ) | ( ~n326 & n335 ) | ( n327 & n335 ) ;
  assign n337 = x30 & n324 ;
  assign n338 = x16 & n337 ;
  assign n339 = ( n94 & ~n101 ) | ( n94 & n338 ) | ( ~n101 & n338 ) ;
  assign n340 = ( n94 & n338 ) | ( n94 & ~n339 ) | ( n338 & ~n339 ) ;
  assign n341 = ( n101 & n339 ) | ( n101 & ~n340 ) | ( n339 & ~n340 ) ;
  assign n342 = ~x32 & n341 ;
  assign n343 = ( x31 & n341 ) | ( x31 & n342 ) | ( n341 & n342 ) ;
  assign n344 = x24 & n324 ;
  assign n345 = x30 & n344 ;
  assign n346 = n123 | n345 ;
  assign n347 = n123 & n345 ;
  assign n348 = n346 & ~n347 ;
  assign n349 = ~x32 & n348 ;
  assign n350 = ( x31 & n348 ) | ( x31 & n349 ) | ( n348 & n349 ) ;
  assign n351 = x26 & n324 ;
  assign n352 = x30 & n351 ;
  assign n353 = n68 | n352 ;
  assign n354 = n68 & n352 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = ~x32 & n355 ;
  assign n357 = ( x31 & n355 ) | ( x31 & n356 ) | ( n355 & n356 ) ;
  assign n358 = x27 & n324 ;
  assign n359 = x30 & n358 ;
  assign n360 = n47 | n359 ;
  assign n361 = n47 & n359 ;
  assign n362 = n360 & ~n361 ;
  assign n363 = ~x32 & n362 ;
  assign n364 = ( x31 & n362 ) | ( x31 & n363 ) | ( n362 & n363 ) ;
  assign n365 = x18 & n337 ;
  assign n366 = ~n165 & n365 ;
  assign n367 = ~x31 & x32 ;
  assign n368 = ( n165 & ~n365 ) | ( n165 & n367 ) | ( ~n365 & n367 ) ;
  assign n369 = ( n366 & ~n367 ) | ( n366 & n368 ) | ( ~n367 & n368 ) ;
  assign n370 = ~x20 & x32 ;
  assign n371 = ( ~x28 & x32 ) | ( ~x28 & n370 ) | ( x32 & n370 ) ;
  assign n372 = n222 | n232 ;
  assign n373 = ( n226 & ~n238 ) | ( n226 & n372 ) | ( ~n238 & n372 ) ;
  assign n374 = n238 | n373 ;
  assign n375 = n186 | n374 ;
  assign n376 = ( ~n193 & n304 ) | ( ~n193 & n375 ) | ( n304 & n375 ) ;
  assign n377 = n193 | n376 ;
  assign n378 = n94 | n377 ;
  assign n379 = ( x32 & n94 ) | ( x32 & ~n377 ) | ( n94 & ~n377 ) ;
  assign n380 = x28 | n94 ;
  assign n381 = ( x32 & n94 ) | ( x32 & n380 ) | ( n94 & n380 ) ;
  assign n382 = ( n378 & n379 ) | ( n378 & ~n381 ) | ( n379 & ~n381 ) ;
  assign n383 = n371 | n382 ;
  assign n384 = n371 & ~n382 ;
  assign n385 = ( ~n371 & n383 ) | ( ~n371 & n384 ) | ( n383 & n384 ) ;
  assign n386 = ~x21 & x32 ;
  assign n387 = ( ~x29 & x32 ) | ( ~x29 & n386 ) | ( x32 & n386 ) ;
  assign n388 = n251 & n300 ;
  assign n389 = ( n251 & n313 ) | ( n251 & n388 ) | ( n313 & n388 ) ;
  assign n390 = n209 | n300 ;
  assign n391 = ( n201 & n209 ) | ( n201 & n390 ) | ( n209 & n390 ) ;
  assign n392 = n263 | n391 ;
  assign n393 = n312 | n392 ;
  assign n394 = n316 | n393 ;
  assign n395 = n389 | n394 ;
  assign n396 = ( ~x8 & x13 ) | ( ~x8 & n135 ) | ( x13 & n135 ) ;
  assign n397 = ( x8 & ~n135 ) | ( x8 & n396 ) | ( ~n135 & n396 ) ;
  assign n398 = ( ~x13 & n396 ) | ( ~x13 & n397 ) | ( n396 & n397 ) ;
  assign n399 = n395 | n398 ;
  assign n400 = ( x32 & ~n395 ) | ( x32 & n398 ) | ( ~n395 & n398 ) ;
  assign n401 = x29 | n398 ;
  assign n402 = ( x32 & n398 ) | ( x32 & n401 ) | ( n398 & n401 ) ;
  assign n403 = ( n399 & n400 ) | ( n399 & ~n402 ) | ( n400 & ~n402 ) ;
  assign n404 = n387 | n403 ;
  assign n405 = n387 & ~n403 ;
  assign n406 = ( ~n387 & n404 ) | ( ~n387 & n405 ) | ( n404 & n405 ) ;
  assign n407 = x25 & n324 ;
  assign n408 = x30 & n407 ;
  assign n409 = n141 & ~n408 ;
  assign n410 = ~n141 & n408 ;
  assign n411 = n409 | n410 ;
  assign n412 = n145 & ~n411 ;
  assign n413 = ( ~n145 & n367 ) | ( ~n145 & n411 ) | ( n367 & n411 ) ;
  assign n414 = ( ~n367 & n412 ) | ( ~n367 & n413 ) | ( n412 & n413 ) ;
  assign y0 = n176 ;
  assign y1 = n184 ;
  assign y2 = n189 ;
  assign y3 = n196 ;
  assign y4 = n206 ;
  assign y5 = n212 ;
  assign y6 = n216 ;
  assign y7 = n225 ;
  assign y8 = n229 ;
  assign y9 = n235 ;
  assign y10 = n241 ;
  assign y11 = n247 ;
  assign y12 = n256 ;
  assign y13 = n260 ;
  assign y14 = n266 ;
  assign y15 = n272 ;
  assign y16 = ~n336 ;
  assign y17 = n343 ;
  assign y18 = n350 ;
  assign y19 = n357 ;
  assign y20 = n364 ;
  assign y21 = n369 ;
  assign y22 = ~n385 ;
  assign y23 = ~n406 ;
  assign y24 = n414 ;
endmodule
