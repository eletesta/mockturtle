module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 ;
  assign n10 = x7 & ~x8 ;
  assign n11 = ~x5 & n10 ;
  assign n12 = ~x3 & n11 ;
  assign n13 = ( x2 & ~x4 ) | ( x2 & n12 ) | ( ~x4 & n12 ) ;
  assign n14 = ~x2 & n13 ;
  assign n15 = x1 | x2 ;
  assign n16 = x3 | n15 ;
  assign n17 = x0 & n16 ;
  assign n18 = x0 | n16 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = x7 | x8 ;
  assign n21 = ( ~x7 & n10 ) | ( ~x7 & n20 ) | ( n10 & n20 ) ;
  assign n22 = ~x4 & x5 ;
  assign n23 = ~x3 & n22 ;
  assign n24 = ~x0 & n23 ;
  assign n25 = ~n15 & n24 ;
  assign n26 = ~x3 & x4 ;
  assign n27 = ~x2 & n26 ;
  assign n28 = ~x0 & n27 ;
  assign n29 = ~x1 & n28 ;
  assign n30 = ( n21 & n25 ) | ( n21 & n29 ) | ( n25 & n29 ) ;
  assign n31 = ~n19 & n30 ;
  assign n32 = ( n19 & n21 ) | ( n19 & n31 ) | ( n21 & n31 ) ;
  assign n33 = ( x0 & x1 ) | ( x0 & ~n32 ) | ( x1 & ~n32 ) ;
  assign n34 = n14 & n33 ;
  assign n35 = ( n14 & n32 ) | ( n14 & ~n34 ) | ( n32 & ~n34 ) ;
  assign n36 = x2 & x3 ;
  assign n37 = ~x3 & x5 ;
  assign n38 = x5 | x8 ;
  assign n39 = x2 & n38 ;
  assign n40 = ( n36 & n37 ) | ( n36 & ~n39 ) | ( n37 & ~n39 ) ;
  assign n41 = x1 | x7 ;
  assign n42 = ( x4 & n40 ) | ( x4 & n41 ) | ( n40 & n41 ) ;
  assign n43 = n40 & ~n42 ;
  assign n44 = ( x2 & ~x5 ) | ( x2 & x7 ) | ( ~x5 & x7 ) ;
  assign n45 = ( ~x4 & x7 ) | ( ~x4 & n44 ) | ( x7 & n44 ) ;
  assign n46 = x7 & ~n45 ;
  assign n47 = n45 | n46 ;
  assign n48 = ( ~x7 & n46 ) | ( ~x7 & n47 ) | ( n46 & n47 ) ;
  assign n49 = ~x6 & x8 ;
  assign n50 = ( x1 & ~n48 ) | ( x1 & n49 ) | ( ~n48 & n49 ) ;
  assign n51 = n48 & n50 ;
  assign n52 = ~x5 & x6 ;
  assign n53 = x2 | x4 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = ( x1 & ~n20 ) | ( x1 & n54 ) | ( ~n20 & n54 ) ;
  assign n56 = ~x1 & n55 ;
  assign n57 = ~x1 & x2 ;
  assign n58 = x6 | n20 ;
  assign n59 = x5 & ~n58 ;
  assign n60 = x3 & ~x4 ;
  assign n61 = n59 & n60 ;
  assign n62 = n57 & n61 ;
  assign n63 = ( ~n51 & n56 ) | ( ~n51 & n62 ) | ( n56 & n62 ) ;
  assign n64 = x3 & ~n62 ;
  assign n65 = ( n51 & n63 ) | ( n51 & ~n64 ) | ( n63 & ~n64 ) ;
  assign n66 = x2 | x3 ;
  assign n67 = x4 & ~x5 ;
  assign n68 = x7 & x8 ;
  assign n69 = x1 & n68 ;
  assign n70 = ( n66 & n67 ) | ( n66 & n69 ) | ( n67 & n69 ) ;
  assign n71 = ~n66 & n70 ;
  assign n72 = ( x1 & x2 ) | ( x1 & ~x7 ) | ( x2 & ~x7 ) ;
  assign n73 = x7 | n72 ;
  assign n74 = ~x1 & x3 ;
  assign n75 = ( ~x2 & n72 ) | ( ~x2 & n74 ) | ( n72 & n74 ) ;
  assign n76 = ( ~x1 & n73 ) | ( ~x1 & n75 ) | ( n73 & n75 ) ;
  assign n77 = x8 & n76 ;
  assign n78 = ( x2 & x3 ) | ( x2 & ~x7 ) | ( x3 & ~x7 ) ;
  assign n79 = ( x2 & x3 ) | ( x2 & x8 ) | ( x3 & x8 ) ;
  assign n80 = n78 & ~n79 ;
  assign n81 = n77 | n80 ;
  assign n82 = ( ~x1 & n77 ) | ( ~x1 & n81 ) | ( n77 & n81 ) ;
  assign n83 = x4 & ~x7 ;
  assign n84 = x1 & x7 ;
  assign n85 = ~x4 & x8 ;
  assign n86 = x1 & ~n85 ;
  assign n87 = ( n83 & n84 ) | ( n83 & ~n86 ) | ( n84 & ~n86 ) ;
  assign n88 = ( ~x2 & n82 ) | ( ~x2 & n87 ) | ( n82 & n87 ) ;
  assign n89 = x3 | n88 ;
  assign n90 = ( ~x3 & n82 ) | ( ~x3 & n89 ) | ( n82 & n89 ) ;
  assign n91 = n71 | n90 ;
  assign n92 = ( ~n43 & n65 ) | ( ~n43 & n91 ) | ( n65 & n91 ) ;
  assign n93 = n43 | n92 ;
  assign n94 = ~x0 & n93 ;
  assign n95 = x3 | x4 ;
  assign n96 = n52 & ~n95 ;
  assign n97 = x2 & n26 ;
  assign n98 = x0 & ~x1 ;
  assign n99 = ~n66 & n98 ;
  assign n100 = ( n36 & ~n97 ) | ( n36 & n99 ) | ( ~n97 & n99 ) ;
  assign n101 = ~x0 & x1 ;
  assign n102 = n99 | n101 ;
  assign n103 = ( n97 & n100 ) | ( n97 & n102 ) | ( n100 & n102 ) ;
  assign n104 = ( ~n23 & n96 ) | ( ~n23 & n103 ) | ( n96 & n103 ) ;
  assign n105 = x1 & x2 ;
  assign n106 = ~x0 & n105 ;
  assign n107 = n103 | n106 ;
  assign n108 = ( n23 & n104 ) | ( n23 & n107 ) | ( n104 & n107 ) ;
  assign n109 = n94 | n108 ;
  assign n110 = ( n21 & n94 ) | ( n21 & n109 ) | ( n94 & n109 ) ;
  assign n111 = ( x4 & x5 ) | ( x4 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n112 = ( ~x3 & x6 ) | ( ~x3 & n111 ) | ( x6 & n111 ) ;
  assign n113 = ( x3 & ~x4 ) | ( x3 & n111 ) | ( ~x4 & n111 ) ;
  assign n114 = n112 | n113 ;
  assign n115 = x2 & ~n114 ;
  assign n116 = ( x0 & x1 ) | ( x0 & n115 ) | ( x1 & n115 ) ;
  assign n117 = ~x0 & n116 ;
  assign n118 = x4 & x5 ;
  assign n119 = x3 & n118 ;
  assign n120 = x0 & ~x3 ;
  assign n121 = x1 & ~x3 ;
  assign n122 = ( n101 & n120 ) | ( n101 & ~n121 ) | ( n120 & ~n121 ) ;
  assign n123 = ( n23 & ~n26 ) | ( n23 & n122 ) | ( ~n26 & n122 ) ;
  assign n124 = n101 | n122 ;
  assign n125 = ( n26 & n123 ) | ( n26 & n124 ) | ( n123 & n124 ) ;
  assign n126 = ~x2 & n125 ;
  assign n127 = n106 | n126 ;
  assign n128 = ( n119 & n126 ) | ( n119 & n127 ) | ( n126 & n127 ) ;
  assign n129 = x3 & ~x7 ;
  assign n130 = x5 & ~x7 ;
  assign n131 = ( n37 & n129 ) | ( n37 & ~n130 ) | ( n129 & ~n130 ) ;
  assign n132 = x8 & n131 ;
  assign n133 = x2 & ~n132 ;
  assign n134 = x5 | n20 ;
  assign n135 = x3 & ~n134 ;
  assign n136 = x2 | n135 ;
  assign n137 = ~n133 & n136 ;
  assign n138 = ( ~x4 & x6 ) | ( ~x4 & n137 ) | ( x6 & n137 ) ;
  assign n139 = x6 & n37 ;
  assign n140 = ( x2 & n68 ) | ( x2 & n139 ) | ( n68 & n139 ) ;
  assign n141 = ~x2 & n140 ;
  assign n142 = x4 & n141 ;
  assign n143 = ( n137 & ~n138 ) | ( n137 & n142 ) | ( ~n138 & n142 ) ;
  assign n144 = x2 & ~n95 ;
  assign n145 = ~x7 & x8 ;
  assign n146 = ( n143 & n144 ) | ( n143 & n145 ) | ( n144 & n145 ) ;
  assign n147 = n52 & ~n146 ;
  assign n148 = ( n52 & n143 ) | ( n52 & ~n147 ) | ( n143 & ~n147 ) ;
  assign n149 = x1 & ~n148 ;
  assign n150 = ( x3 & x6 ) | ( x3 & x8 ) | ( x6 & x8 ) ;
  assign n151 = ( ~x7 & x8 ) | ( ~x7 & n150 ) | ( x8 & n150 ) ;
  assign n152 = x8 & ~n151 ;
  assign n153 = n151 | n152 ;
  assign n154 = ( ~x8 & n152 ) | ( ~x8 & n153 ) | ( n152 & n153 ) ;
  assign n155 = x2 & ~x5 ;
  assign n156 = x2 & ~n155 ;
  assign n157 = n154 & n156 ;
  assign n158 = ( x3 & x6 ) | ( x3 & ~x7 ) | ( x6 & ~x7 ) ;
  assign n159 = ~n150 & n158 ;
  assign n160 = ( ~n155 & n156 ) | ( ~n155 & n159 ) | ( n156 & n159 ) ;
  assign n161 = ( ~x5 & n157 ) | ( ~x5 & n160 ) | ( n157 & n160 ) ;
  assign n162 = ~x4 & n161 ;
  assign n163 = x1 | n162 ;
  assign n164 = ~n149 & n163 ;
  assign n165 = ( ~x1 & x5 ) | ( ~x1 & x7 ) | ( x5 & x7 ) ;
  assign n166 = ( x2 & x5 ) | ( x2 & n165 ) | ( x5 & n165 ) ;
  assign n167 = ( x1 & ~x2 ) | ( x1 & n166 ) | ( ~x2 & n166 ) ;
  assign n168 = ~x7 & n167 ;
  assign n169 = ( ~x5 & n166 ) | ( ~x5 & n168 ) | ( n166 & n168 ) ;
  assign n170 = x4 | n169 ;
  assign n171 = ~x5 & x7 ;
  assign n172 = n105 & n171 ;
  assign n173 = x4 & ~n172 ;
  assign n174 = n170 & ~n173 ;
  assign n175 = ( x3 & ~x8 ) | ( x3 & n174 ) | ( ~x8 & n174 ) ;
  assign n176 = x5 & ~n20 ;
  assign n177 = ( x1 & ~n53 ) | ( x1 & n176 ) | ( ~n53 & n176 ) ;
  assign n178 = ~x1 & n177 ;
  assign n179 = ~x3 & n178 ;
  assign n180 = ( n174 & ~n175 ) | ( n174 & n179 ) | ( ~n175 & n179 ) ;
  assign n181 = ( x1 & x4 ) | ( x1 & ~x8 ) | ( x4 & ~x8 ) ;
  assign n182 = ( x2 & x8 ) | ( x2 & n181 ) | ( x8 & n181 ) ;
  assign n183 = ( x1 & x4 ) | ( x1 & n182 ) | ( x4 & n182 ) ;
  assign n184 = n181 & ~n183 ;
  assign n185 = ( n182 & ~n183 ) | ( n182 & n184 ) | ( ~n183 & n184 ) ;
  assign n186 = x3 | n185 ;
  assign n187 = x4 & x8 ;
  assign n188 = ( x2 & x4 ) | ( x2 & n187 ) | ( x4 & n187 ) ;
  assign n189 = ~x1 & n188 ;
  assign n190 = x3 & ~n189 ;
  assign n191 = n186 & ~n190 ;
  assign n192 = x3 & x4 ;
  assign n193 = ( x2 & ~x8 ) | ( x2 & n15 ) | ( ~x8 & n15 ) ;
  assign n194 = ( x2 & x8 ) | ( x2 & ~n15 ) | ( x8 & ~n15 ) ;
  assign n195 = ( ~x2 & n193 ) | ( ~x2 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ( x3 & x4 ) | ( x3 & n195 ) | ( x4 & n195 ) ;
  assign n197 = ( n191 & ~n192 ) | ( n191 & n196 ) | ( ~n192 & n196 ) ;
  assign n198 = x7 | n197 ;
  assign n199 = ( x1 & ~x2 ) | ( x1 & x3 ) | ( ~x2 & x3 ) ;
  assign n200 = x1 & ~n199 ;
  assign n201 = x2 & x4 ;
  assign n202 = ( ~x3 & n199 ) | ( ~x3 & n201 ) | ( n199 & n201 ) ;
  assign n203 = ( x2 & ~n200 ) | ( x2 & n202 ) | ( ~n200 & n202 ) ;
  assign n204 = x8 & ~n203 ;
  assign n205 = x7 & ~n204 ;
  assign n206 = n198 & ~n205 ;
  assign n207 = ( ~x0 & n180 ) | ( ~x0 & n206 ) | ( n180 & n206 ) ;
  assign n208 = ~n164 & n207 ;
  assign n209 = ( ~x0 & n164 ) | ( ~x0 & n208 ) | ( n164 & n208 ) ;
  assign n210 = ( ~n117 & n128 ) | ( ~n117 & n209 ) | ( n128 & n209 ) ;
  assign n211 = n21 | n209 ;
  assign n212 = ( n117 & n210 ) | ( n117 & n211 ) | ( n210 & n211 ) ;
  assign n213 = ( x3 & x5 ) | ( x3 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n214 = x5 & ~n213 ;
  assign n215 = ( ~x7 & x8 ) | ( ~x7 & n214 ) | ( x8 & n214 ) ;
  assign n216 = ( ~n213 & n214 ) | ( ~n213 & n215 ) | ( n214 & n215 ) ;
  assign n217 = x2 & n216 ;
  assign n218 = ( x3 & ~x7 ) | ( x3 & x8 ) | ( ~x7 & x8 ) ;
  assign n219 = ( ~x5 & x8 ) | ( ~x5 & n218 ) | ( x8 & n218 ) ;
  assign n220 = x8 & ~n219 ;
  assign n221 = n219 | n220 ;
  assign n222 = ( ~x8 & n220 ) | ( ~x8 & n221 ) | ( n220 & n221 ) ;
  assign n223 = x2 | n222 ;
  assign n224 = ( ~x2 & n217 ) | ( ~x2 & n223 ) | ( n217 & n223 ) ;
  assign n225 = x1 & ~n224 ;
  assign n226 = x5 & n10 ;
  assign n227 = x2 & ~x3 ;
  assign n228 = n226 & n227 ;
  assign n229 = x1 | n228 ;
  assign n230 = ~n225 & n229 ;
  assign n231 = x4 & ~n230 ;
  assign n232 = ( x3 & x5 ) | ( x3 & x7 ) | ( x5 & x7 ) ;
  assign n233 = ( x3 & x8 ) | ( x3 & ~n232 ) | ( x8 & ~n232 ) ;
  assign n234 = ( ~x7 & x8 ) | ( ~x7 & n232 ) | ( x8 & n232 ) ;
  assign n235 = ~n233 & n234 ;
  assign n236 = x2 & ~n235 ;
  assign n237 = n136 & ~n236 ;
  assign n238 = ~x1 & n237 ;
  assign n239 = x4 | n238 ;
  assign n240 = ~n231 & n239 ;
  assign n241 = x6 & ~n240 ;
  assign n242 = x4 | x7 ;
  assign n243 = ( ~x4 & n83 ) | ( ~x4 & n242 ) | ( n83 & n242 ) ;
  assign n244 = x8 | n243 ;
  assign n245 = x5 | n244 ;
  assign n246 = x2 & n245 ;
  assign n247 = x5 & n68 ;
  assign n248 = x4 & n247 ;
  assign n249 = x2 | n248 ;
  assign n250 = ~n246 & n249 ;
  assign n251 = x3 & n250 ;
  assign n252 = n11 | n251 ;
  assign n253 = ( n144 & n251 ) | ( n144 & n252 ) | ( n251 & n252 ) ;
  assign n254 = x1 & n253 ;
  assign n255 = x6 | n254 ;
  assign n256 = ~n241 & n255 ;
  assign n257 = x0 & n256 ;
  assign n258 = x6 & n10 ;
  assign n259 = n22 & n99 ;
  assign n260 = n258 & n259 ;
  assign n261 = x2 & n60 ;
  assign n262 = x0 & x1 ;
  assign n263 = x1 & ~n262 ;
  assign n264 = n261 & n263 ;
  assign n265 = ( n27 & ~n262 ) | ( n27 & n263 ) | ( ~n262 & n263 ) ;
  assign n266 = ( x0 & n264 ) | ( x0 & n265 ) | ( n264 & n265 ) ;
  assign n267 = ~n21 & n266 ;
  assign n268 = ( x3 & ~x5 ) | ( x3 & x8 ) | ( ~x5 & x8 ) ;
  assign n269 = n218 & ~n268 ;
  assign n270 = ( x3 & x7 ) | ( x3 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n271 = ( x4 & ~x8 ) | ( x4 & n270 ) | ( ~x8 & n270 ) ;
  assign n272 = x8 & n271 ;
  assign n273 = n271 & ~n272 ;
  assign n274 = ( x8 & ~n272 ) | ( x8 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = ( x2 & ~x5 ) | ( x2 & n274 ) | ( ~x5 & n274 ) ;
  assign n276 = x4 & n10 ;
  assign n277 = ~n66 & n276 ;
  assign n278 = ~x5 & n277 ;
  assign n279 = ( ~n274 & n275 ) | ( ~n274 & n278 ) | ( n275 & n278 ) ;
  assign n280 = ( x2 & x4 ) | ( x2 & ~n279 ) | ( x4 & ~n279 ) ;
  assign n281 = n269 & n280 ;
  assign n282 = ( n269 & n279 ) | ( n269 & ~n281 ) | ( n279 & ~n281 ) ;
  assign n283 = ( ~x0 & x1 ) | ( ~x0 & n282 ) | ( x1 & n282 ) ;
  assign n284 = x5 & n145 ;
  assign n285 = ~x2 & x4 ;
  assign n286 = x4 & ~n285 ;
  assign n287 = n284 & n286 ;
  assign n288 = ( n11 & ~n285 ) | ( n11 & n286 ) | ( ~n285 & n286 ) ;
  assign n289 = ( ~x2 & n287 ) | ( ~x2 & n288 ) | ( n287 & n288 ) ;
  assign n290 = x3 | n289 ;
  assign n291 = ( x4 & x7 ) | ( x4 & x8 ) | ( x7 & x8 ) ;
  assign n292 = ( x5 & ~x8 ) | ( x5 & n291 ) | ( ~x8 & n291 ) ;
  assign n293 = ( x4 & x7 ) | ( x4 & n292 ) | ( x7 & n292 ) ;
  assign n294 = ~n291 & n293 ;
  assign n295 = ( ~n292 & n293 ) | ( ~n292 & n294 ) | ( n293 & n294 ) ;
  assign n296 = ~x2 & n295 ;
  assign n297 = x3 & ~n296 ;
  assign n298 = n290 & ~n297 ;
  assign n299 = ( x0 & x1 ) | ( x0 & ~n298 ) | ( x1 & ~n298 ) ;
  assign n300 = n283 & ~n299 ;
  assign n301 = ( x3 & x8 ) | ( x3 & n242 ) | ( x8 & n242 ) ;
  assign n302 = x7 & ~n301 ;
  assign n303 = ( ~x4 & n242 ) | ( ~x4 & n301 ) | ( n242 & n301 ) ;
  assign n304 = ( ~x7 & n302 ) | ( ~x7 & n303 ) | ( n302 & n303 ) ;
  assign n305 = ( ~x1 & x2 ) | ( ~x1 & n304 ) | ( x2 & n304 ) ;
  assign n306 = ~x3 & x8 ;
  assign n307 = ( ~x4 & x7 ) | ( ~x4 & n306 ) | ( x7 & n306 ) ;
  assign n308 = ( x4 & ~x8 ) | ( x4 & n306 ) | ( ~x8 & n306 ) ;
  assign n309 = ( x3 & n307 ) | ( x3 & n308 ) | ( n307 & n308 ) ;
  assign n310 = ( x1 & x2 ) | ( x1 & ~n309 ) | ( x2 & ~n309 ) ;
  assign n311 = n305 & ~n310 ;
  assign n312 = x2 | x8 ;
  assign n313 = ( x4 & ~x7 ) | ( x4 & n312 ) | ( ~x7 & n312 ) ;
  assign n314 = ( x2 & x4 ) | ( x2 & ~n312 ) | ( x4 & ~n312 ) ;
  assign n315 = ( x8 & ~n313 ) | ( x8 & n314 ) | ( ~n313 & n314 ) ;
  assign n316 = ( x1 & ~x3 ) | ( x1 & n315 ) | ( ~x3 & n315 ) ;
  assign n317 = ( ~x2 & n20 ) | ( ~x2 & n53 ) | ( n20 & n53 ) ;
  assign n318 = ( x1 & x3 ) | ( x1 & ~n317 ) | ( x3 & ~n317 ) ;
  assign n319 = n316 & n318 ;
  assign n320 = x0 & ~n15 ;
  assign n321 = ~n95 & n320 ;
  assign n322 = n145 & n321 ;
  assign n323 = ( ~n311 & n319 ) | ( ~n311 & n322 ) | ( n319 & n322 ) ;
  assign n324 = x0 & ~n322 ;
  assign n325 = ( n311 & n323 ) | ( n311 & ~n324 ) | ( n323 & ~n324 ) ;
  assign n326 = n300 | n325 ;
  assign n327 = ( n266 & ~n267 ) | ( n266 & n326 ) | ( ~n267 & n326 ) ;
  assign n328 = n260 | n327 ;
  assign n329 = ( n256 & ~n257 ) | ( n256 & n328 ) | ( ~n257 & n328 ) ;
  assign n330 = x4 & ~x6 ;
  assign n331 = ~x5 & n68 ;
  assign n332 = ( ~x3 & x5 ) | ( ~x3 & x8 ) | ( x5 & x8 ) ;
  assign n333 = ( x4 & ~x8 ) | ( x4 & n332 ) | ( ~x8 & n332 ) ;
  assign n334 = ( x4 & x5 ) | ( x4 & ~n332 ) | ( x5 & ~n332 ) ;
  assign n335 = n333 & ~n334 ;
  assign n336 = ( ~x1 & x7 ) | ( ~x1 & n335 ) | ( x7 & n335 ) ;
  assign n337 = x4 & n74 ;
  assign n338 = ( x5 & x8 ) | ( x5 & n337 ) | ( x8 & n337 ) ;
  assign n339 = ~x8 & n338 ;
  assign n340 = ~x7 & n339 ;
  assign n341 = ( n335 & ~n336 ) | ( n335 & n340 ) | ( ~n336 & n340 ) ;
  assign n342 = ( ~x1 & n60 ) | ( ~x1 & n341 ) | ( n60 & n341 ) ;
  assign n343 = n331 & ~n342 ;
  assign n344 = ( n331 & n341 ) | ( n331 & ~n343 ) | ( n341 & ~n343 ) ;
  assign n345 = x2 & ~n344 ;
  assign n346 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n347 = ( x3 & x4 ) | ( x3 & ~x8 ) | ( x4 & ~x8 ) ;
  assign n348 = n346 & ~n347 ;
  assign n349 = x5 & n348 ;
  assign n350 = ~x1 & n349 ;
  assign n351 = x2 | n350 ;
  assign n352 = ~n345 & n351 ;
  assign n353 = ( ~x0 & x6 ) | ( ~x0 & n352 ) | ( x6 & n352 ) ;
  assign n354 = ~x1 & x4 ;
  assign n355 = x4 & ~n354 ;
  assign n356 = n131 & n355 ;
  assign n357 = x5 | x7 ;
  assign n358 = ( n354 & ~n355 ) | ( n354 & n357 ) | ( ~n355 & n357 ) ;
  assign n359 = ( x1 & ~n356 ) | ( x1 & n358 ) | ( ~n356 & n358 ) ;
  assign n360 = ~x2 & n359 ;
  assign n361 = ( x1 & x3 ) | ( x1 & x5 ) | ( x3 & x5 ) ;
  assign n362 = ( ~x3 & x7 ) | ( ~x3 & n361 ) | ( x7 & n361 ) ;
  assign n363 = ( x1 & x5 ) | ( x1 & n362 ) | ( x5 & n362 ) ;
  assign n364 = n361 & ~n363 ;
  assign n365 = ( n362 & ~n363 ) | ( n362 & n364 ) | ( ~n363 & n364 ) ;
  assign n366 = ~x4 & n365 ;
  assign n367 = x2 & ~n366 ;
  assign n368 = n360 | n367 ;
  assign n369 = x8 | n368 ;
  assign n370 = ~x3 & n247 ;
  assign n371 = ~x4 & n370 ;
  assign n372 = n369 & ~n371 ;
  assign n373 = ( x1 & n369 ) | ( x1 & n372 ) | ( n369 & n372 ) ;
  assign n374 = ( x0 & x6 ) | ( x0 & n373 ) | ( x6 & n373 ) ;
  assign n375 = n353 & ~n374 ;
  assign n376 = x3 | x5 ;
  assign n377 = x4 | n376 ;
  assign n378 = x0 & x2 ;
  assign n379 = x0 & ~n378 ;
  assign n380 = ~n377 & n379 ;
  assign n381 = ( n119 & ~n378 ) | ( n119 & n379 ) | ( ~n378 & n379 ) ;
  assign n382 = ( x2 & n380 ) | ( x2 & n381 ) | ( n380 & n381 ) ;
  assign n383 = x1 | n382 ;
  assign n384 = ( x2 & x4 ) | ( x2 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n385 = x5 | n384 ;
  assign n386 = ( x2 & x3 ) | ( x2 & ~n385 ) | ( x3 & ~n385 ) ;
  assign n387 = ( n384 & n385 ) | ( n384 & ~n386 ) | ( n385 & ~n386 ) ;
  assign n388 = x0 | n387 ;
  assign n389 = x1 & n388 ;
  assign n390 = n383 & ~n389 ;
  assign n391 = ~x7 & n390 ;
  assign n392 = n106 & ~n357 ;
  assign n393 = ~n95 & n392 ;
  assign n394 = x4 & x7 ;
  assign n395 = ( x4 & x8 ) | ( x4 & ~n285 ) | ( x8 & ~n285 ) ;
  assign n396 = ( x7 & ~x8 ) | ( x7 & n285 ) | ( ~x8 & n285 ) ;
  assign n397 = ( ~n394 & n395 ) | ( ~n394 & n396 ) | ( n395 & n396 ) ;
  assign n398 = x5 & n397 ;
  assign n399 = ( ~x2 & x7 ) | ( ~x2 & x8 ) | ( x7 & x8 ) ;
  assign n400 = ~x7 & n399 ;
  assign n401 = ( x2 & n399 ) | ( x2 & n400 ) | ( n399 & n400 ) ;
  assign n402 = x4 & n401 ;
  assign n403 = x5 | n402 ;
  assign n404 = ~n398 & n403 ;
  assign n405 = ( n22 & n83 ) | ( n22 & ~n130 ) | ( n83 & ~n130 ) ;
  assign n406 = ( x2 & x8 ) | ( x2 & n405 ) | ( x8 & n405 ) ;
  assign n407 = ( x0 & ~x8 ) | ( x0 & n406 ) | ( ~x8 & n406 ) ;
  assign n408 = ( x0 & x2 ) | ( x0 & ~n406 ) | ( x2 & ~n406 ) ;
  assign n409 = n407 & ~n408 ;
  assign n410 = x0 & ~n409 ;
  assign n411 = ( n404 & n409 ) | ( n404 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = x3 | n411 ;
  assign n413 = x8 & n53 ;
  assign n414 = ( n68 & n83 ) | ( n68 & ~n413 ) | ( n83 & ~n413 ) ;
  assign n415 = x5 | n414 ;
  assign n416 = n20 | n53 ;
  assign n417 = x5 & n416 ;
  assign n418 = n415 & ~n417 ;
  assign n419 = ~x0 & n418 ;
  assign n420 = x3 & ~n419 ;
  assign n421 = n412 & ~n420 ;
  assign n422 = x1 | n421 ;
  assign n423 = n144 & ~n284 ;
  assign n424 = ( ~x2 & x4 ) | ( ~x2 & x5 ) | ( x4 & x5 ) ;
  assign n425 = ( x2 & ~x7 ) | ( x2 & n424 ) | ( ~x7 & n424 ) ;
  assign n426 = ( x4 & x5 ) | ( x4 & n425 ) | ( x5 & n425 ) ;
  assign n427 = ~n424 & n426 ;
  assign n428 = ( ~n425 & n426 ) | ( ~n425 & n427 ) | ( n426 & n427 ) ;
  assign n429 = ( ~x3 & x8 ) | ( ~x3 & n428 ) | ( x8 & n428 ) ;
  assign n430 = x4 & ~n66 ;
  assign n431 = ~n357 & n430 ;
  assign n432 = ~x8 & n431 ;
  assign n433 = ( n428 & ~n429 ) | ( n428 & n432 ) | ( ~n429 & n432 ) ;
  assign n434 = x2 & ~n201 ;
  assign n435 = n331 & n434 ;
  assign n436 = ( n176 & ~n201 ) | ( n176 & n434 ) | ( ~n201 & n434 ) ;
  assign n437 = ( x4 & n435 ) | ( x4 & n436 ) | ( n435 & n436 ) ;
  assign n438 = n433 | n437 ;
  assign n439 = ( n144 & ~n423 ) | ( n144 & n438 ) | ( ~n423 & n438 ) ;
  assign n440 = ~x0 & n439 ;
  assign n441 = x1 & ~n440 ;
  assign n442 = n422 & ~n441 ;
  assign n443 = n393 | n442 ;
  assign n444 = ( n390 & ~n391 ) | ( n390 & n443 ) | ( ~n391 & n443 ) ;
  assign n445 = x4 | x6 ;
  assign n446 = ( ~x4 & n330 ) | ( ~x4 & n445 ) | ( n330 & n445 ) ;
  assign n447 = ~x2 & x8 ;
  assign n448 = ( x3 & n446 ) | ( x3 & ~n447 ) | ( n446 & ~n447 ) ;
  assign n449 = n446 & ~n448 ;
  assign n450 = x1 | n449 ;
  assign n451 = x6 | x8 ;
  assign n452 = x4 & ~n451 ;
  assign n453 = n36 & n452 ;
  assign n454 = x1 & ~n453 ;
  assign n455 = n450 & ~n454 ;
  assign n456 = ( ~x5 & n130 ) | ( ~x5 & n357 ) | ( n130 & n357 ) ;
  assign n457 = ( x0 & n455 ) | ( x0 & ~n456 ) | ( n455 & ~n456 ) ;
  assign n458 = x8 & n26 ;
  assign n459 = ( x6 & n320 ) | ( x6 & n458 ) | ( n320 & n458 ) ;
  assign n460 = ~x6 & n459 ;
  assign n461 = n456 & n460 ;
  assign n462 = ( n455 & ~n457 ) | ( n455 & n461 ) | ( ~n457 & n461 ) ;
  assign n463 = ~x4 & x6 ;
  assign n464 = n145 & n463 ;
  assign n465 = ( x1 & x2 ) | ( x1 & ~x8 ) | ( x2 & ~x8 ) ;
  assign n466 = n72 & ~n465 ;
  assign n467 = ( n10 & ~n15 ) | ( n10 & n466 ) | ( ~n15 & n466 ) ;
  assign n468 = x3 & ~n467 ;
  assign n469 = ( x3 & n466 ) | ( x3 & ~n468 ) | ( n466 & ~n468 ) ;
  assign n470 = x4 & x6 ;
  assign n471 = x6 & ~n470 ;
  assign n472 = n469 & n471 ;
  assign n473 = ( x2 & x3 ) | ( x2 & ~x8 ) | ( x3 & ~x8 ) ;
  assign n474 = ~x3 & n473 ;
  assign n475 = ( x1 & x2 ) | ( x1 & ~n474 ) | ( x2 & ~n474 ) ;
  assign n476 = ( n473 & n474 ) | ( n473 & ~n475 ) | ( n474 & ~n475 ) ;
  assign n477 = x7 | n466 ;
  assign n478 = ( n466 & n476 ) | ( n466 & n477 ) | ( n476 & n477 ) ;
  assign n479 = ( ~n470 & n471 ) | ( ~n470 & n478 ) | ( n471 & n478 ) ;
  assign n480 = ( x4 & n472 ) | ( x4 & n479 ) | ( n472 & n479 ) ;
  assign n481 = ~x0 & n480 ;
  assign n482 = n99 | n481 ;
  assign n483 = ( n464 & n481 ) | ( n464 & n482 ) | ( n481 & n482 ) ;
  assign n484 = n462 | n483 ;
  assign n485 = ( ~n375 & n444 ) | ( ~n375 & n484 ) | ( n444 & n484 ) ;
  assign n486 = n375 | n485 ;
  assign n487 = ( x2 & x7 ) | ( x2 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n488 = ( x5 & x7 ) | ( x5 & x8 ) | ( x7 & x8 ) ;
  assign n489 = ~n487 & n488 ;
  assign n490 = ( x2 & x5 ) | ( x2 & n21 ) | ( x5 & n21 ) ;
  assign n491 = ( x0 & ~x5 ) | ( x0 & n490 ) | ( ~x5 & n490 ) ;
  assign n492 = ( x0 & x2 ) | ( x0 & ~n490 ) | ( x2 & ~n490 ) ;
  assign n493 = n491 & ~n492 ;
  assign n494 = x0 & ~n493 ;
  assign n495 = ( n489 & n493 ) | ( n489 & ~n494 ) | ( n493 & ~n494 ) ;
  assign n496 = x1 | n495 ;
  assign n497 = ( x5 & x7 ) | ( x5 & ~n399 ) | ( x7 & ~n399 ) ;
  assign n498 = ( ~x7 & x8 ) | ( ~x7 & n497 ) | ( x8 & n497 ) ;
  assign n499 = n399 & n498 ;
  assign n500 = x5 & ~n499 ;
  assign n501 = ( n497 & n499 ) | ( n497 & ~n500 ) | ( n499 & ~n500 ) ;
  assign n502 = ~x0 & n501 ;
  assign n503 = x1 & ~n502 ;
  assign n504 = n496 & ~n503 ;
  assign n505 = x3 | n504 ;
  assign n506 = ( x1 & x2 ) | ( x1 & x8 ) | ( x2 & x8 ) ;
  assign n507 = ( x7 & ~x8 ) | ( x7 & n506 ) | ( ~x8 & n506 ) ;
  assign n508 = ( x1 & x2 ) | ( x1 & n507 ) | ( x2 & n507 ) ;
  assign n509 = n506 & ~n508 ;
  assign n510 = ( n507 & ~n508 ) | ( n507 & n509 ) | ( ~n508 & n509 ) ;
  assign n511 = x1 & ~x2 ;
  assign n512 = n510 | n511 ;
  assign n513 = ( n247 & n510 ) | ( n247 & n512 ) | ( n510 & n512 ) ;
  assign n514 = ~x0 & n513 ;
  assign n515 = x3 & ~n514 ;
  assign n516 = n505 & ~n515 ;
  assign n517 = ( x4 & ~x6 ) | ( x4 & n516 ) | ( ~x6 & n516 ) ;
  assign n518 = ( ~n330 & n486 ) | ( ~n330 & n517 ) | ( n486 & n517 ) ;
  assign n519 = ( x0 & ~x4 ) | ( x0 & x5 ) | ( ~x4 & x5 ) ;
  assign n520 = ( ~x3 & x5 ) | ( ~x3 & n519 ) | ( x5 & n519 ) ;
  assign n521 = x5 & ~n520 ;
  assign n522 = n520 | n521 ;
  assign n523 = ( ~x5 & n521 ) | ( ~x5 & n522 ) | ( n521 & n522 ) ;
  assign n524 = x2 | n523 ;
  assign n525 = ( x3 & ~x4 ) | ( x3 & x5 ) | ( ~x4 & x5 ) ;
  assign n526 = x6 | n525 ;
  assign n527 = ( ~x5 & x6 ) | ( ~x5 & n525 ) | ( x6 & n525 ) ;
  assign n528 = ( x5 & ~n526 ) | ( x5 & n527 ) | ( ~n526 & n527 ) ;
  assign n529 = ~x0 & n528 ;
  assign n530 = x2 & ~n529 ;
  assign n531 = n524 & ~n530 ;
  assign n532 = x1 | n531 ;
  assign n533 = ( ~x2 & x3 ) | ( ~x2 & x5 ) | ( x3 & x5 ) ;
  assign n534 = ( x2 & ~x4 ) | ( x2 & n533 ) | ( ~x4 & n533 ) ;
  assign n535 = ( x3 & x5 ) | ( x3 & n534 ) | ( x5 & n534 ) ;
  assign n536 = ~n533 & n535 ;
  assign n537 = ( ~n534 & n535 ) | ( ~n534 & n536 ) | ( n535 & n536 ) ;
  assign n538 = x6 & ~n537 ;
  assign n539 = x2 & ~x4 ;
  assign n540 = ( x4 & ~n26 ) | ( x4 & n539 ) | ( ~n26 & n539 ) ;
  assign n541 = x5 | n540 ;
  assign n542 = ~x6 & n541 ;
  assign n543 = n538 | n542 ;
  assign n544 = x0 | n543 ;
  assign n545 = x1 & n544 ;
  assign n546 = n532 & ~n545 ;
  assign n547 = n21 & n546 ;
  assign n548 = ~x6 & n456 ;
  assign n549 = x4 & ~n201 ;
  assign n550 = n548 & n549 ;
  assign n551 = ~x6 & x7 ;
  assign n552 = ~x5 & n551 ;
  assign n553 = x6 & n130 ;
  assign n554 = n552 | n553 ;
  assign n555 = ( ~n201 & n549 ) | ( ~n201 & n554 ) | ( n549 & n554 ) ;
  assign n556 = ( x2 & n550 ) | ( x2 & n555 ) | ( n550 & n555 ) ;
  assign n557 = x1 & ~n556 ;
  assign n558 = ( x4 & x5 ) | ( x4 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n559 = x4 & ~n558 ;
  assign n560 = ( x5 & x6 ) | ( x5 & n559 ) | ( x6 & n559 ) ;
  assign n561 = ( ~n558 & n559 ) | ( ~n558 & n560 ) | ( n559 & n560 ) ;
  assign n562 = ~x2 & n561 ;
  assign n563 = x1 | n562 ;
  assign n564 = ~n557 & n563 ;
  assign n565 = ( x0 & ~x3 ) | ( x0 & n564 ) | ( ~x3 & n564 ) ;
  assign n566 = x6 | x7 ;
  assign n567 = ~n66 & n67 ;
  assign n568 = ( x1 & ~n566 ) | ( x1 & n567 ) | ( ~n566 & n567 ) ;
  assign n569 = ~x1 & n568 ;
  assign n570 = ~x0 & n569 ;
  assign n571 = ( n564 & ~n565 ) | ( n564 & n570 ) | ( ~n565 & n570 ) ;
  assign n572 = x6 & x7 ;
  assign n573 = n99 & n572 ;
  assign n574 = n67 & n573 ;
  assign n575 = x6 & n145 ;
  assign n576 = ~x1 & x5 ;
  assign n577 = ( n74 & n227 ) | ( n74 & ~n576 ) | ( n227 & ~n576 ) ;
  assign n578 = ( ~x2 & n227 ) | ( ~x2 & n577 ) | ( n227 & n577 ) ;
  assign n579 = ~x4 & n578 ;
  assign n580 = ~x0 & n579 ;
  assign n581 = ( ~x3 & n118 ) | ( ~x3 & n580 ) | ( n118 & n580 ) ;
  assign n582 = n320 & ~n581 ;
  assign n583 = ( n320 & n580 ) | ( n320 & ~n582 ) | ( n580 & ~n582 ) ;
  assign n584 = ~x6 & n10 ;
  assign n585 = n583 & n584 ;
  assign n586 = ( n575 & n583 ) | ( n575 & n585 ) | ( n583 & n585 ) ;
  assign n587 = x5 | x6 ;
  assign n588 = ( x2 & x6 ) | ( x2 & x8 ) | ( x6 & x8 ) ;
  assign n589 = x5 & x8 ;
  assign n590 = ( ~x6 & n588 ) | ( ~x6 & n589 ) | ( n588 & n589 ) ;
  assign n591 = ( ~x2 & x6 ) | ( ~x2 & x7 ) | ( x6 & x7 ) ;
  assign n592 = x2 & n591 ;
  assign n593 = ( x5 & x6 ) | ( x5 & ~n592 ) | ( x6 & ~n592 ) ;
  assign n594 = ( n591 & n592 ) | ( n591 & ~n593 ) | ( n592 & ~n593 ) ;
  assign n595 = ( x4 & ~x8 ) | ( x4 & n594 ) | ( ~x8 & n594 ) ;
  assign n596 = x5 & x6 ;
  assign n597 = x6 & ~x7 ;
  assign n598 = ( ~x2 & n596 ) | ( ~x2 & n597 ) | ( n596 & n597 ) ;
  assign n599 = ( ~x2 & x7 ) | ( ~x2 & n596 ) | ( x7 & n596 ) ;
  assign n600 = ( x7 & n598 ) | ( x7 & ~n599 ) | ( n598 & ~n599 ) ;
  assign n601 = ( x4 & x8 ) | ( x4 & ~n600 ) | ( x8 & ~n600 ) ;
  assign n602 = n595 & ~n601 ;
  assign n603 = ( x4 & x7 ) | ( x4 & ~n602 ) | ( x7 & ~n602 ) ;
  assign n604 = n590 & n603 ;
  assign n605 = ( n590 & n602 ) | ( n590 & ~n604 ) | ( n602 & ~n604 ) ;
  assign n606 = ( ~x0 & x3 ) | ( ~x0 & n605 ) | ( x3 & n605 ) ;
  assign n607 = ( x5 & ~x7 ) | ( x5 & x8 ) | ( ~x7 & x8 ) ;
  assign n608 = ( x2 & x7 ) | ( x2 & n607 ) | ( x7 & n607 ) ;
  assign n609 = ( x7 & x8 ) | ( x7 & ~n608 ) | ( x8 & ~n608 ) ;
  assign n610 = n607 & n609 ;
  assign n611 = ( x2 & ~n608 ) | ( x2 & n610 ) | ( ~n608 & n610 ) ;
  assign n612 = x6 | n611 ;
  assign n613 = x5 & ~x8 ;
  assign n614 = ( ~x5 & n38 ) | ( ~x5 & n613 ) | ( n38 & n613 ) ;
  assign n615 = x7 & n614 ;
  assign n616 = x2 & n615 ;
  assign n617 = x6 & ~n616 ;
  assign n618 = n612 & ~n617 ;
  assign n619 = x4 | n618 ;
  assign n620 = ( x5 & x6 ) | ( x5 & ~x8 ) | ( x6 & ~x8 ) ;
  assign n621 = ( x2 & ~x5 ) | ( x2 & n620 ) | ( ~x5 & n620 ) ;
  assign n622 = ( x5 & x8 ) | ( x5 & n621 ) | ( x8 & n621 ) ;
  assign n623 = n620 & ~n622 ;
  assign n624 = ( x2 & ~n621 ) | ( x2 & n623 ) | ( ~n621 & n623 ) ;
  assign n625 = x7 & n624 ;
  assign n626 = x4 & ~n625 ;
  assign n627 = n619 & ~n626 ;
  assign n628 = ( x0 & x3 ) | ( x0 & ~n627 ) | ( x3 & ~n627 ) ;
  assign n629 = n606 & ~n628 ;
  assign n630 = x2 | n95 ;
  assign n631 = x0 & ~n630 ;
  assign n632 = ( n145 & n629 ) | ( n145 & n631 ) | ( n629 & n631 ) ;
  assign n633 = n587 | n632 ;
  assign n634 = ( ~n587 & n629 ) | ( ~n587 & n633 ) | ( n629 & n633 ) ;
  assign n635 = x1 | n634 ;
  assign n636 = ( x4 & ~x5 ) | ( x4 & x6 ) | ( ~x5 & x6 ) ;
  assign n637 = ( x5 & ~x7 ) | ( x5 & n636 ) | ( ~x7 & n636 ) ;
  assign n638 = ( x4 & x6 ) | ( x4 & n637 ) | ( x6 & n637 ) ;
  assign n639 = n636 & ~n638 ;
  assign n640 = ( n637 & ~n638 ) | ( n637 & n639 ) | ( ~n638 & n639 ) ;
  assign n641 = x3 & n640 ;
  assign n642 = ( x4 & x5 ) | ( x4 & x6 ) | ( x5 & x6 ) ;
  assign n643 = ( x4 & ~x7 ) | ( x4 & n596 ) | ( ~x7 & n596 ) ;
  assign n644 = n642 & ~n643 ;
  assign n645 = x3 | n644 ;
  assign n646 = ( ~x3 & n641 ) | ( ~x3 & n645 ) | ( n641 & n645 ) ;
  assign n647 = x8 | n646 ;
  assign n648 = ( x6 & x7 ) | ( x6 & ~n642 ) | ( x7 & ~n642 ) ;
  assign n649 = ( x4 & x5 ) | ( x4 & ~n648 ) | ( x5 & ~n648 ) ;
  assign n650 = ~n642 & n649 ;
  assign n651 = ( n648 & n649 ) | ( n648 & n650 ) | ( n649 & n650 ) ;
  assign n652 = ~x3 & n651 ;
  assign n653 = x8 & ~n652 ;
  assign n654 = n647 & ~n653 ;
  assign n655 = x2 & n192 ;
  assign n656 = n11 & ~n630 ;
  assign n657 = n284 | n656 ;
  assign n658 = ( n655 & n656 ) | ( n655 & n657 ) | ( n656 & n657 ) ;
  assign n659 = ( x2 & n654 ) | ( x2 & n658 ) | ( n654 & n658 ) ;
  assign n660 = ( ~x3 & x4 ) | ( ~x3 & x6 ) | ( x4 & x6 ) ;
  assign n661 = ( x4 & x7 ) | ( x4 & ~n660 ) | ( x7 & ~n660 ) ;
  assign n662 = ( x3 & ~x6 ) | ( x3 & n661 ) | ( ~x6 & n661 ) ;
  assign n663 = n660 & n662 ;
  assign n664 = ( ~n661 & n662 ) | ( ~n661 & n663 ) | ( n662 & n663 ) ;
  assign n665 = x8 | n664 ;
  assign n666 = ( x3 & x7 ) | ( x3 & n60 ) | ( x7 & n60 ) ;
  assign n667 = ( ~x3 & x7 ) | ( ~x3 & n60 ) | ( x7 & n60 ) ;
  assign n668 = ( x3 & ~n666 ) | ( x3 & n667 ) | ( ~n666 & n667 ) ;
  assign n669 = x6 & n668 ;
  assign n670 = x8 & ~n669 ;
  assign n671 = n665 & ~n670 ;
  assign n672 = x3 & ~x5 ;
  assign n673 = ( x4 & n584 ) | ( x4 & n672 ) | ( n584 & n672 ) ;
  assign n674 = ~x4 & n673 ;
  assign n675 = x5 | n674 ;
  assign n676 = ( n671 & n674 ) | ( n671 & n675 ) | ( n674 & n675 ) ;
  assign n677 = ( ~x2 & n658 ) | ( ~x2 & n676 ) | ( n658 & n676 ) ;
  assign n678 = n659 | n677 ;
  assign n679 = ~x0 & n678 ;
  assign n680 = x1 & ~n679 ;
  assign n681 = n635 & ~n680 ;
  assign n682 = n586 | n681 ;
  assign n683 = ( ~n571 & n574 ) | ( ~n571 & n682 ) | ( n574 & n682 ) ;
  assign n684 = n571 | n683 ;
  assign n685 = ( x2 & x6 ) | ( x2 & ~x8 ) | ( x6 & ~x8 ) ;
  assign n686 = ( ~x2 & x4 ) | ( ~x2 & n685 ) | ( x4 & n685 ) ;
  assign n687 = ( ~x4 & x8 ) | ( ~x4 & n685 ) | ( x8 & n685 ) ;
  assign n688 = n686 & n687 ;
  assign n689 = x4 & ~x8 ;
  assign n690 = ( x0 & x2 ) | ( x0 & n689 ) | ( x2 & n689 ) ;
  assign n691 = ( x2 & x4 ) | ( x2 & ~n690 ) | ( x4 & ~n690 ) ;
  assign n692 = ( x0 & ~x8 ) | ( x0 & n691 ) | ( ~x8 & n691 ) ;
  assign n693 = ~n690 & n692 ;
  assign n694 = ( ~x5 & x6 ) | ( ~x5 & n693 ) | ( x6 & n693 ) ;
  assign n695 = ~x5 & x8 ;
  assign n696 = x4 & n695 ;
  assign n697 = ( x0 & x2 ) | ( x0 & n696 ) | ( x2 & n696 ) ;
  assign n698 = ~x0 & n697 ;
  assign n699 = ~x6 & n698 ;
  assign n700 = ( n693 & ~n694 ) | ( n693 & n699 ) | ( ~n694 & n699 ) ;
  assign n701 = ( x0 & x5 ) | ( x0 & ~n700 ) | ( x5 & ~n700 ) ;
  assign n702 = n688 & n701 ;
  assign n703 = ( n688 & n700 ) | ( n688 & ~n702 ) | ( n700 & ~n702 ) ;
  assign n704 = x3 | n703 ;
  assign n705 = ( ~x2 & x5 ) | ( ~x2 & x6 ) | ( x5 & x6 ) ;
  assign n706 = ( x2 & x4 ) | ( x2 & n705 ) | ( x4 & n705 ) ;
  assign n707 = ( x5 & x6 ) | ( x5 & n706 ) | ( x6 & n706 ) ;
  assign n708 = n705 & ~n707 ;
  assign n709 = ( n706 & ~n707 ) | ( n706 & n708 ) | ( ~n707 & n708 ) ;
  assign n710 = ~x8 & n709 ;
  assign n711 = ~x0 & n710 ;
  assign n712 = x3 & ~n711 ;
  assign n713 = n704 & ~n712 ;
  assign n714 = x1 | n713 ;
  assign n715 = x2 & ~x8 ;
  assign n716 = x2 & ~n715 ;
  assign n717 = x4 & n716 ;
  assign n718 = ( x6 & ~n715 ) | ( x6 & n716 ) | ( ~n715 & n716 ) ;
  assign n719 = ( ~x8 & n717 ) | ( ~x8 & n718 ) | ( n717 & n718 ) ;
  assign n720 = x3 & n719 ;
  assign n721 = ( x2 & x4 ) | ( x2 & x8 ) | ( x4 & x8 ) ;
  assign n722 = ( x4 & ~x6 ) | ( x4 & n721 ) | ( ~x6 & n721 ) ;
  assign n723 = x4 & ~n722 ;
  assign n724 = n722 | n723 ;
  assign n725 = ( ~x4 & n723 ) | ( ~x4 & n724 ) | ( n723 & n724 ) ;
  assign n726 = x3 | n725 ;
  assign n727 = ( ~x3 & n720 ) | ( ~x3 & n726 ) | ( n720 & n726 ) ;
  assign n728 = x5 | n727 ;
  assign n729 = x6 & ~x8 ;
  assign n730 = n655 & n729 ;
  assign n731 = x5 & ~n730 ;
  assign n732 = n728 & ~n731 ;
  assign n733 = ~x0 & n732 ;
  assign n734 = x1 & ~n733 ;
  assign n735 = n714 & ~n734 ;
  assign n736 = n684 | n735 ;
  assign n737 = ( n546 & ~n547 ) | ( n546 & n736 ) | ( ~n547 & n736 ) ;
  assign n738 = x5 & x7 ;
  assign n739 = ( ~x5 & n26 ) | ( ~x5 & n738 ) | ( n26 & n738 ) ;
  assign n740 = ~x1 & n739 ;
  assign n741 = ~x2 & n740 ;
  assign n742 = x0 & n741 ;
  assign n743 = ( ~x1 & x2 ) | ( ~x1 & x7 ) | ( x2 & x7 ) ;
  assign n744 = ~x2 & n743 ;
  assign n745 = ( x1 & ~x5 ) | ( x1 & n744 ) | ( ~x5 & n744 ) ;
  assign n746 = ( n743 & n744 ) | ( n743 & n745 ) | ( n744 & n745 ) ;
  assign n747 = ( ~x3 & x4 ) | ( ~x3 & n746 ) | ( x4 & n746 ) ;
  assign n748 = ( x1 & ~x2 ) | ( x1 & x5 ) | ( ~x2 & x5 ) ;
  assign n749 = n44 & ~n748 ;
  assign n750 = x7 & ~n749 ;
  assign n751 = ( n748 & n749 ) | ( n748 & ~n750 ) | ( n749 & ~n750 ) ;
  assign n752 = ( x3 & x4 ) | ( x3 & n751 ) | ( x4 & n751 ) ;
  assign n753 = n747 & ~n752 ;
  assign n754 = ( ~n118 & n130 ) | ( ~n118 & n242 ) | ( n130 & n242 ) ;
  assign n755 = ( x2 & x3 ) | ( x2 & ~n754 ) | ( x3 & ~n754 ) ;
  assign n756 = ( x1 & ~x3 ) | ( x1 & n755 ) | ( ~x3 & n755 ) ;
  assign n757 = ( x1 & x2 ) | ( x1 & ~n755 ) | ( x2 & ~n755 ) ;
  assign n758 = n756 & ~n757 ;
  assign n759 = n753 | n758 ;
  assign n760 = ~x0 & n759 ;
  assign n761 = n742 | n760 ;
  assign n762 = ( ~x6 & n451 ) | ( ~x6 & n729 ) | ( n451 & n729 ) ;
  assign n763 = n761 & n762 ;
  assign n764 = x4 | x5 ;
  assign n765 = ( x2 & x3 ) | ( x2 & n764 ) | ( x3 & n764 ) ;
  assign n766 = ( x2 & x3 ) | ( x2 & ~n764 ) | ( x3 & ~n764 ) ;
  assign n767 = ( x4 & x5 ) | ( x4 & n766 ) | ( x5 & n766 ) ;
  assign n768 = n765 & ~n767 ;
  assign n769 = x1 & n768 ;
  assign n770 = x2 | x5 ;
  assign n771 = ( x2 & n60 ) | ( x2 & ~n770 ) | ( n60 & ~n770 ) ;
  assign n772 = x1 | n771 ;
  assign n773 = ( ~x1 & n769 ) | ( ~x1 & n772 ) | ( n769 & n772 ) ;
  assign n774 = ( ~x0 & x7 ) | ( ~x0 & n773 ) | ( x7 & n773 ) ;
  assign n775 = x2 | n37 ;
  assign n776 = ( x2 & ~x4 ) | ( x2 & n37 ) | ( ~x4 & n37 ) ;
  assign n777 = n775 & ~n776 ;
  assign n778 = ( ~x2 & n775 ) | ( ~x2 & n777 ) | ( n775 & n777 ) ;
  assign n779 = x1 | n778 ;
  assign n780 = x2 & n119 ;
  assign n781 = x1 & ~n780 ;
  assign n782 = n779 & ~n781 ;
  assign n783 = ( x0 & x7 ) | ( x0 & ~n782 ) | ( x7 & ~n782 ) ;
  assign n784 = n774 & ~n783 ;
  assign n785 = ~x4 & x7 ;
  assign n786 = x2 & x5 ;
  assign n787 = ( x3 & ~n101 ) | ( x3 & n786 ) | ( ~n101 & n786 ) ;
  assign n788 = n101 & n787 ;
  assign n789 = ~x3 & n98 ;
  assign n790 = ( x2 & ~x5 ) | ( x2 & n789 ) | ( ~x5 & n789 ) ;
  assign n791 = ~x2 & n790 ;
  assign n792 = n788 | n791 ;
  assign n793 = ( ~x4 & x7 ) | ( ~x4 & n792 ) | ( x7 & n792 ) ;
  assign n794 = ( n785 & n792 ) | ( n785 & ~n793 ) | ( n792 & ~n793 ) ;
  assign n795 = n784 | n794 ;
  assign n796 = ( ~x6 & x8 ) | ( ~x6 & n795 ) | ( x8 & n795 ) ;
  assign n797 = ( n49 & n795 ) | ( n49 & ~n796 ) | ( n795 & ~n796 ) ;
  assign n798 = ( x2 & x3 ) | ( x2 & x7 ) | ( x3 & x7 ) ;
  assign n799 = ( ~x5 & x7 ) | ( ~x5 & n798 ) | ( x7 & n798 ) ;
  assign n800 = x7 & ~n799 ;
  assign n801 = n799 | n800 ;
  assign n802 = ( ~x7 & n800 ) | ( ~x7 & n801 ) | ( n800 & n801 ) ;
  assign n803 = ( x1 & x6 ) | ( x1 & ~n802 ) | ( x6 & ~n802 ) ;
  assign n804 = x3 & n57 ;
  assign n805 = ~n357 & n804 ;
  assign n806 = x6 & n805 ;
  assign n807 = ( n802 & n803 ) | ( n802 & n806 ) | ( n803 & n806 ) ;
  assign n808 = x3 | n587 ;
  assign n809 = ( x1 & x2 ) | ( x1 & ~n808 ) | ( x2 & ~n808 ) ;
  assign n810 = ~x1 & n809 ;
  assign n811 = x5 & ~n566 ;
  assign n812 = ~x2 & x5 ;
  assign n813 = ( ~x3 & x4 ) | ( ~x3 & n812 ) | ( x4 & n812 ) ;
  assign n814 = ( x2 & x3 ) | ( x2 & n813 ) | ( x3 & n813 ) ;
  assign n815 = ( x4 & x5 ) | ( x4 & ~n814 ) | ( x5 & ~n814 ) ;
  assign n816 = ~n813 & n815 ;
  assign n817 = x4 & n227 ;
  assign n818 = n171 & n817 ;
  assign n819 = x7 & ~n818 ;
  assign n820 = ( n816 & n818 ) | ( n816 & ~n819 ) | ( n818 & ~n819 ) ;
  assign n821 = x6 & n820 ;
  assign n822 = n261 | n821 ;
  assign n823 = ( n811 & n821 ) | ( n811 & n822 ) | ( n821 & n822 ) ;
  assign n824 = x8 & n823 ;
  assign n825 = x5 & ~x6 ;
  assign n826 = ( ~n22 & n463 ) | ( ~n22 & n825 ) | ( n463 & n825 ) ;
  assign n827 = ( ~x2 & x7 ) | ( ~x2 & n826 ) | ( x7 & n826 ) ;
  assign n828 = ~x7 & n827 ;
  assign n829 = ( x2 & x3 ) | ( x2 & n828 ) | ( x3 & n828 ) ;
  assign n830 = ( n827 & n828 ) | ( n827 & n829 ) | ( n828 & n829 ) ;
  assign n831 = ( x2 & ~x5 ) | ( x2 & n26 ) | ( ~x5 & n26 ) ;
  assign n832 = ( x2 & x3 ) | ( x2 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n833 = ( ~x3 & x4 ) | ( ~x3 & n831 ) | ( x4 & n831 ) ;
  assign n834 = ( n26 & n832 ) | ( n26 & ~n833 ) | ( n832 & ~n833 ) ;
  assign n835 = n831 & ~n834 ;
  assign n836 = ( ~x6 & n830 ) | ( ~x6 & n835 ) | ( n830 & n835 ) ;
  assign n837 = x7 | n836 ;
  assign n838 = ( ~x7 & n830 ) | ( ~x7 & n837 ) | ( n830 & n837 ) ;
  assign n839 = x8 | n838 ;
  assign n840 = ( ~x8 & n824 ) | ( ~x8 & n839 ) | ( n824 & n839 ) ;
  assign n841 = x1 & n840 ;
  assign n842 = ~x2 & x3 ;
  assign n843 = ( x2 & x7 ) | ( x2 & n812 ) | ( x7 & n812 ) ;
  assign n844 = ( x3 & x7 ) | ( x3 & n812 ) | ( x7 & n812 ) ;
  assign n845 = ( n842 & n843 ) | ( n842 & ~n844 ) | ( n843 & ~n844 ) ;
  assign n846 = ~n66 & n552 ;
  assign n847 = x6 | n846 ;
  assign n848 = ( n845 & n846 ) | ( n845 & n847 ) | ( n846 & n847 ) ;
  assign n849 = ( x4 & ~x8 ) | ( x4 & n848 ) | ( ~x8 & n848 ) ;
  assign n850 = x2 & ~n58 ;
  assign n851 = n37 & n850 ;
  assign n852 = ~x4 & n851 ;
  assign n853 = ( n848 & ~n849 ) | ( n848 & n852 ) | ( ~n849 & n852 ) ;
  assign n854 = ( x5 & x6 ) | ( x5 & ~n607 ) | ( x6 & ~n607 ) ;
  assign n855 = ( x7 & ~x8 ) | ( x7 & n854 ) | ( ~x8 & n854 ) ;
  assign n856 = n607 & n855 ;
  assign n857 = ( ~n854 & n855 ) | ( ~n854 & n856 ) | ( n855 & n856 ) ;
  assign n858 = x2 & n857 ;
  assign n859 = ( ~x6 & x7 ) | ( ~x6 & x8 ) | ( x7 & x8 ) ;
  assign n860 = ( x5 & x6 ) | ( x5 & ~n859 ) | ( x6 & ~n859 ) ;
  assign n861 = ( ~x6 & n695 ) | ( ~x6 & n860 ) | ( n695 & n860 ) ;
  assign n862 = x2 | n861 ;
  assign n863 = ( ~x2 & n858 ) | ( ~x2 & n862 ) | ( n858 & n862 ) ;
  assign n864 = ( ~x3 & x4 ) | ( ~x3 & n863 ) | ( x4 & n863 ) ;
  assign n865 = ( x6 & ~x7 ) | ( x6 & x8 ) | ( ~x7 & x8 ) ;
  assign n866 = ( x2 & ~x8 ) | ( x2 & n865 ) | ( ~x8 & n865 ) ;
  assign n867 = ( x2 & x6 ) | ( x2 & ~n865 ) | ( x6 & ~n865 ) ;
  assign n868 = n866 & ~n867 ;
  assign n869 = x5 & ~n868 ;
  assign n870 = ~x2 & n68 ;
  assign n871 = x5 | n870 ;
  assign n872 = ~n869 & n871 ;
  assign n873 = ( x3 & x4 ) | ( x3 & n872 ) | ( x4 & n872 ) ;
  assign n874 = n864 & n873 ;
  assign n875 = n853 | n874 ;
  assign n876 = ~x1 & n875 ;
  assign n877 = n841 | n876 ;
  assign n878 = ( ~n807 & n810 ) | ( ~n807 & n877 ) | ( n810 & n877 ) ;
  assign n879 = x4 | x8 ;
  assign n880 = ( ~x4 & n689 ) | ( ~x4 & n879 ) | ( n689 & n879 ) ;
  assign n881 = n877 | n880 ;
  assign n882 = ( n807 & n878 ) | ( n807 & n881 ) | ( n878 & n881 ) ;
  assign n883 = x0 & n882 ;
  assign n884 = ~x6 & n68 ;
  assign n885 = n259 & n884 ;
  assign n886 = x0 & x5 ;
  assign n887 = ( x3 & ~x6 ) | ( x3 & n886 ) | ( ~x6 & n886 ) ;
  assign n888 = ( x0 & x3 ) | ( x0 & ~n887 ) | ( x3 & ~n887 ) ;
  assign n889 = ( x5 & ~x6 ) | ( x5 & n888 ) | ( ~x6 & n888 ) ;
  assign n890 = ~n887 & n889 ;
  assign n891 = ~x7 & n890 ;
  assign n892 = x1 | n891 ;
  assign n893 = ( x3 & ~n376 ) | ( x3 & n572 ) | ( ~n376 & n572 ) ;
  assign n894 = ~x0 & n893 ;
  assign n895 = x1 & ~n894 ;
  assign n896 = n892 & ~n895 ;
  assign n897 = x2 | n896 ;
  assign n898 = ( x1 & x5 ) | ( x1 & x6 ) | ( x5 & x6 ) ;
  assign n899 = ( ~x1 & x3 ) | ( ~x1 & n898 ) | ( x3 & n898 ) ;
  assign n900 = ( x5 & x6 ) | ( x5 & n899 ) | ( x6 & n899 ) ;
  assign n901 = ~n898 & n900 ;
  assign n902 = ( ~n899 & n900 ) | ( ~n899 & n901 ) | ( n900 & n901 ) ;
  assign n903 = x7 & n902 ;
  assign n904 = ~x0 & n903 ;
  assign n905 = x2 & ~n904 ;
  assign n906 = n897 & ~n905 ;
  assign n907 = ~x4 & n906 ;
  assign n908 = ( x2 & x6 ) | ( x2 & ~x7 ) | ( x6 & ~x7 ) ;
  assign n909 = ( x2 & ~x5 ) | ( x2 & x6 ) | ( ~x5 & x6 ) ;
  assign n910 = ~n908 & n909 ;
  assign n911 = x1 & x4 ;
  assign n912 = ( x3 & ~n910 ) | ( x3 & n911 ) | ( ~n910 & n911 ) ;
  assign n913 = n910 & n912 ;
  assign n914 = n907 | n913 ;
  assign n915 = ( ~x0 & n907 ) | ( ~x0 & n914 ) | ( n907 & n914 ) ;
  assign n916 = n885 | n915 ;
  assign n917 = ( n882 & ~n883 ) | ( n882 & n916 ) | ( ~n883 & n916 ) ;
  assign n918 = n797 | n917 ;
  assign n919 = ( n761 & ~n763 ) | ( n761 & n918 ) | ( ~n763 & n918 ) ;
  assign n920 = x6 & x8 ;
  assign n921 = x1 & ~x4 ;
  assign n922 = x3 & n921 ;
  assign n923 = ( ~x1 & x2 ) | ( ~x1 & n921 ) | ( x2 & n921 ) ;
  assign n924 = ( ~x3 & n511 ) | ( ~x3 & n923 ) | ( n511 & n923 ) ;
  assign n925 = ( x3 & ~n922 ) | ( x3 & n924 ) | ( ~n922 & n924 ) ;
  assign n926 = ( x1 & x2 ) | ( x1 & ~x4 ) | ( x2 & ~x4 ) ;
  assign n927 = ( x1 & ~x5 ) | ( x1 & n926 ) | ( ~x5 & n926 ) ;
  assign n928 = x1 & ~n927 ;
  assign n929 = n927 | n928 ;
  assign n930 = ( ~x1 & n928 ) | ( ~x1 & n929 ) | ( n928 & n929 ) ;
  assign n931 = x5 & ~n930 ;
  assign n932 = ( n925 & ~n930 ) | ( n925 & n931 ) | ( ~n930 & n931 ) ;
  assign n933 = x8 & ~n932 ;
  assign n934 = ( n26 & ~n155 ) | ( n26 & n766 ) | ( ~n155 & n766 ) ;
  assign n935 = x1 | n934 ;
  assign n936 = x3 & n22 ;
  assign n937 = x2 & n936 ;
  assign n938 = x1 & ~n937 ;
  assign n939 = n935 & ~n938 ;
  assign n940 = x8 | n939 ;
  assign n941 = ( ~x8 & n933 ) | ( ~x8 & n940 ) | ( n933 & n940 ) ;
  assign n942 = ( ~x0 & x6 ) | ( ~x0 & n941 ) | ( x6 & n941 ) ;
  assign n943 = ( ~x2 & x3 ) | ( ~x2 & x8 ) | ( x3 & x8 ) ;
  assign n944 = n533 & ~n943 ;
  assign n945 = ( x2 & x3 ) | ( x2 & ~n36 ) | ( x3 & ~n36 ) ;
  assign n946 = ( x1 & ~x4 ) | ( x1 & n945 ) | ( ~x4 & n945 ) ;
  assign n947 = ~n36 & n946 ;
  assign n948 = ( ~x5 & x8 ) | ( ~x5 & n947 ) | ( x8 & n947 ) ;
  assign n949 = ( x1 & x3 ) | ( x1 & x4 ) | ( x3 & x4 ) ;
  assign n950 = ( ~x2 & x4 ) | ( ~x2 & n949 ) | ( x4 & n949 ) ;
  assign n951 = x4 & ~n950 ;
  assign n952 = n950 | n951 ;
  assign n953 = ( ~x4 & n951 ) | ( ~x4 & n952 ) | ( n951 & n952 ) ;
  assign n954 = ( x5 & x8 ) | ( x5 & n953 ) | ( x8 & n953 ) ;
  assign n955 = n948 & n954 ;
  assign n956 = ( x1 & ~x4 ) | ( x1 & n955 ) | ( ~x4 & n955 ) ;
  assign n957 = n944 & ~n956 ;
  assign n958 = ( n944 & n955 ) | ( n944 & ~n957 ) | ( n955 & ~n957 ) ;
  assign n959 = ( x0 & x6 ) | ( x0 & ~n958 ) | ( x6 & ~n958 ) ;
  assign n960 = n942 & ~n959 ;
  assign n961 = ~x4 & n306 ;
  assign n962 = ( x1 & ~x4 ) | ( x1 & x8 ) | ( ~x4 & x8 ) ;
  assign n963 = x8 & ~n962 ;
  assign n964 = ( x1 & x2 ) | ( x1 & n963 ) | ( x2 & n963 ) ;
  assign n965 = ( ~n962 & n963 ) | ( ~n962 & n964 ) | ( n963 & n964 ) ;
  assign n966 = x3 & n965 ;
  assign n967 = ~x0 & n966 ;
  assign n968 = n15 & ~n967 ;
  assign n969 = ( n961 & n967 ) | ( n961 & ~n968 ) | ( n967 & ~n968 ) ;
  assign n970 = ( x5 & x6 ) | ( x5 & ~n969 ) | ( x6 & ~n969 ) ;
  assign n971 = ( n587 & n960 ) | ( n587 & ~n970 ) | ( n960 & ~n970 ) ;
  assign n972 = x7 & ~n971 ;
  assign n973 = ( ~x4 & x5 ) | ( ~x4 & x6 ) | ( x5 & x6 ) ;
  assign n974 = x4 & n973 ;
  assign n975 = ( x3 & ~x6 ) | ( x3 & n974 ) | ( ~x6 & n974 ) ;
  assign n976 = ( n973 & n974 ) | ( n973 & n975 ) | ( n974 & n975 ) ;
  assign n977 = ~x2 & n976 ;
  assign n978 = ( x4 & x5 ) | ( x4 & ~x8 ) | ( x5 & ~x8 ) ;
  assign n979 = ( ~x5 & x6 ) | ( ~x5 & x8 ) | ( x6 & x8 ) ;
  assign n980 = ~x4 & n979 ;
  assign n981 = n978 | n980 ;
  assign n982 = ( x2 & x3 ) | ( x2 & ~n981 ) | ( x3 & ~n981 ) ;
  assign n983 = x5 | n451 ;
  assign n984 = x4 & ~n983 ;
  assign n985 = x2 & n984 ;
  assign n986 = ~x3 & n985 ;
  assign n987 = ( n981 & n982 ) | ( n981 & ~n986 ) | ( n982 & ~n986 ) ;
  assign n988 = ~x4 & n842 ;
  assign n989 = ~n587 & n988 ;
  assign n990 = n987 & ~n989 ;
  assign n991 = ( ~n976 & n977 ) | ( ~n976 & n990 ) | ( n977 & n990 ) ;
  assign n992 = x1 & ~n991 ;
  assign n993 = ( ~x6 & n285 ) | ( ~x6 & n614 ) | ( n285 & n614 ) ;
  assign n994 = ~n614 & n993 ;
  assign n995 = ( n539 & n920 ) | ( n539 & n994 ) | ( n920 & n994 ) ;
  assign n996 = x5 & ~n995 ;
  assign n997 = ( x5 & n994 ) | ( x5 & ~n996 ) | ( n994 & ~n996 ) ;
  assign n998 = ( x4 & x6 ) | ( x4 & x8 ) | ( x6 & x8 ) ;
  assign n999 = x8 & n998 ;
  assign n1000 = ( x2 & x4 ) | ( x2 & n998 ) | ( x4 & n998 ) ;
  assign n1001 = x8 | n1000 ;
  assign n1002 = ~n999 & n1001 ;
  assign n1003 = x3 | n1002 ;
  assign n1004 = x2 & n187 ;
  assign n1005 = x3 & ~n1004 ;
  assign n1006 = n1003 & ~n1005 ;
  assign n1007 = x5 | n1006 ;
  assign n1008 = ~n630 & n920 ;
  assign n1009 = x5 & ~n1008 ;
  assign n1010 = n1007 & ~n1009 ;
  assign n1011 = n997 | n1010 ;
  assign n1012 = ~x1 & n1011 ;
  assign n1013 = n992 | n1012 ;
  assign n1014 = ~x0 & n1013 ;
  assign n1015 = x7 | n1014 ;
  assign n1016 = ~n972 & n1015 ;
  assign n1017 = ( x0 & x4 ) | ( x0 & x5 ) | ( x4 & x5 ) ;
  assign n1018 = ( x4 & x7 ) | ( x4 & ~n1017 ) | ( x7 & ~n1017 ) ;
  assign n1019 = ( x0 & x5 ) | ( x0 & ~n1018 ) | ( x5 & ~n1018 ) ;
  assign n1020 = ~n1017 & n1019 ;
  assign n1021 = ( n1018 & n1019 ) | ( n1018 & n1020 ) | ( n1019 & n1020 ) ;
  assign n1022 = x1 & n1021 ;
  assign n1023 = ( x0 & x4 ) | ( x0 & n456 ) | ( x4 & n456 ) ;
  assign n1024 = ( x1 & ~x4 ) | ( x1 & n1023 ) | ( ~x4 & n1023 ) ;
  assign n1025 = ( x0 & x1 ) | ( x0 & ~n1023 ) | ( x1 & ~n1023 ) ;
  assign n1026 = n1024 & ~n1025 ;
  assign n1027 = ~x4 & n101 ;
  assign n1028 = ~n357 & n1027 ;
  assign n1029 = n1026 | n1028 ;
  assign n1030 = ( n1021 & ~n1022 ) | ( n1021 & n1029 ) | ( ~n1022 & n1029 ) ;
  assign n1031 = x2 | n1030 ;
  assign n1032 = ( x1 & x5 ) | ( x1 & ~n394 ) | ( x5 & ~n394 ) ;
  assign n1033 = ( x1 & ~x5 ) | ( x1 & x7 ) | ( ~x5 & x7 ) ;
  assign n1034 = x1 & ~n1033 ;
  assign n1035 = n1032 & ~n1034 ;
  assign n1036 = ~x0 & n1035 ;
  assign n1037 = x2 & ~n1036 ;
  assign n1038 = n1031 & ~n1037 ;
  assign n1039 = x3 | n1038 ;
  assign n1040 = x5 & n785 ;
  assign n1041 = ~x2 & n1040 ;
  assign n1042 = ( ~x2 & n67 ) | ( ~x2 & n1041 ) | ( n67 & n1041 ) ;
  assign n1043 = x1 & ~n1042 ;
  assign n1044 = ( x2 & x5 ) | ( x2 & x7 ) | ( x5 & x7 ) ;
  assign n1045 = x4 & n1044 ;
  assign n1046 = ( n53 & n738 ) | ( n53 & ~n1045 ) | ( n738 & ~n1045 ) ;
  assign n1047 = x1 | n1046 ;
  assign n1048 = ( ~x1 & n1043 ) | ( ~x1 & n1047 ) | ( n1043 & n1047 ) ;
  assign n1049 = x0 | n1048 ;
  assign n1050 = x3 & n1049 ;
  assign n1051 = n1039 & ~n1050 ;
  assign n1052 = ( x6 & x8 ) | ( x6 & n1051 ) | ( x8 & n1051 ) ;
  assign n1053 = ( ~n920 & n1016 ) | ( ~n920 & n1052 ) | ( n1016 & n1052 ) ;
  assign n1054 = ( ~x1 & x2 ) | ( ~x1 & x5 ) | ( x2 & x5 ) ;
  assign n1055 = ( x5 & x7 ) | ( x5 & ~n1054 ) | ( x7 & ~n1054 ) ;
  assign n1056 = ( ~x2 & x7 ) | ( ~x2 & n1054 ) | ( x7 & n1054 ) ;
  assign n1057 = n1055 & ~n1056 ;
  assign n1058 = x0 & n1057 ;
  assign n1059 = x7 & n98 ;
  assign n1060 = ( x2 & x5 ) | ( x2 & n1059 ) | ( x5 & n1059 ) ;
  assign n1061 = ~x2 & n1060 ;
  assign n1062 = ( x0 & x1 ) | ( x0 & x4 ) | ( x1 & x4 ) ;
  assign n1063 = ( x0 & x7 ) | ( x0 & ~n1062 ) | ( x7 & ~n1062 ) ;
  assign n1064 = ( ~x1 & x7 ) | ( ~x1 & n1062 ) | ( x7 & n1062 ) ;
  assign n1065 = ~n1063 & n1064 ;
  assign n1066 = ( x0 & x1 ) | ( x0 & ~n1065 ) | ( x1 & ~n1065 ) ;
  assign n1067 = n1040 & n1066 ;
  assign n1068 = ( n1040 & n1065 ) | ( n1040 & ~n1067 ) | ( n1065 & ~n1067 ) ;
  assign n1069 = x2 | n1068 ;
  assign n1070 = ( x1 & x4 ) | ( x1 & ~x7 ) | ( x4 & ~x7 ) ;
  assign n1071 = ( ~x4 & x5 ) | ( ~x4 & n1070 ) | ( x5 & n1070 ) ;
  assign n1072 = ( x1 & x5 ) | ( x1 & ~n1070 ) | ( x5 & ~n1070 ) ;
  assign n1073 = n1071 & ~n1072 ;
  assign n1074 = ~x0 & n1073 ;
  assign n1075 = x2 & ~n1074 ;
  assign n1076 = n1069 & ~n1075 ;
  assign n1077 = n1061 | n1076 ;
  assign n1078 = ( n1057 & ~n1058 ) | ( n1057 & n1077 ) | ( ~n1058 & n1077 ) ;
  assign n1079 = x3 | n1078 ;
  assign n1080 = x2 & ~x7 ;
  assign n1081 = ( ~x2 & n67 ) | ( ~x2 & n1080 ) | ( n67 & n1080 ) ;
  assign n1082 = x1 & n1081 ;
  assign n1083 = ( x2 & ~x4 ) | ( x2 & x7 ) | ( ~x4 & x7 ) ;
  assign n1084 = ( x5 & ~x7 ) | ( x5 & n1083 ) | ( ~x7 & n1083 ) ;
  assign n1085 = ( x2 & ~x4 ) | ( x2 & n1084 ) | ( ~x4 & n1084 ) ;
  assign n1086 = ~n1083 & n1085 ;
  assign n1087 = ( ~n1084 & n1085 ) | ( ~n1084 & n1086 ) | ( n1085 & n1086 ) ;
  assign n1088 = x1 | n1087 ;
  assign n1089 = ( ~x1 & n1082 ) | ( ~x1 & n1088 ) | ( n1082 & n1088 ) ;
  assign n1090 = ~x0 & n1089 ;
  assign n1091 = x3 & ~n1090 ;
  assign n1092 = n1079 & ~n1091 ;
  assign n1093 = n1053 | n1092 ;
  assign n1094 = ( ~n762 & n1053 ) | ( ~n762 & n1093 ) | ( n1053 & n1093 ) ;
  assign n1095 = x0 & ~x6 ;
  assign n1096 = ( ~x4 & x7 ) | ( ~x4 & n1095 ) | ( x7 & n1095 ) ;
  assign n1097 = ( x6 & ~x7 ) | ( x6 & n1095 ) | ( ~x7 & n1095 ) ;
  assign n1098 = ( ~x0 & x4 ) | ( ~x0 & n1097 ) | ( x4 & n1097 ) ;
  assign n1099 = n1096 | n1098 ;
  assign n1100 = ~x3 & n1099 ;
  assign n1101 = ~x4 & n551 ;
  assign n1102 = ~x0 & n1101 ;
  assign n1103 = x3 & ~n1102 ;
  assign n1104 = n1100 | n1103 ;
  assign n1105 = ~x2 & n1104 ;
  assign n1106 = ( x3 & x4 ) | ( x3 & ~x7 ) | ( x4 & ~x7 ) ;
  assign n1107 = ( ~x3 & x6 ) | ( ~x3 & n1106 ) | ( x6 & n1106 ) ;
  assign n1108 = ( ~x6 & x7 ) | ( ~x6 & n1106 ) | ( x7 & n1106 ) ;
  assign n1109 = n1107 & n1108 ;
  assign n1110 = ~x0 & n1109 ;
  assign n1111 = x2 & ~n1110 ;
  assign n1112 = n1105 | n1111 ;
  assign n1113 = ~x1 & n1112 ;
  assign n1114 = x4 & n129 ;
  assign n1115 = x2 & ~n1114 ;
  assign n1116 = ~x4 & n572 ;
  assign n1117 = ~x3 & n1116 ;
  assign n1118 = x2 | n1117 ;
  assign n1119 = ~n1115 & n1118 ;
  assign n1120 = ~x0 & n1119 ;
  assign n1121 = x1 & ~n1120 ;
  assign n1122 = n1113 | n1121 ;
  assign n1123 = n614 | n1122 ;
  assign n1124 = ( ~x0 & x5 ) | ( ~x0 & x7 ) | ( x5 & x7 ) ;
  assign n1125 = ( x7 & x8 ) | ( x7 & ~n1124 ) | ( x8 & ~n1124 ) ;
  assign n1126 = ( x0 & ~x5 ) | ( x0 & n1125 ) | ( ~x5 & n1125 ) ;
  assign n1127 = n1124 & n1126 ;
  assign n1128 = ( ~n1125 & n1126 ) | ( ~n1125 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = ~x4 & n1128 ;
  assign n1130 = x1 | n1129 ;
  assign n1131 = x7 & ~n614 ;
  assign n1132 = x4 & n1131 ;
  assign n1133 = ~x0 & n1132 ;
  assign n1134 = x1 & ~n1133 ;
  assign n1135 = n1130 & ~n1134 ;
  assign n1136 = x3 | n1135 ;
  assign n1137 = x1 & ~n67 ;
  assign n1138 = ( n67 & n68 ) | ( n67 & n1137 ) | ( n68 & n1137 ) ;
  assign n1139 = ~x0 & n1138 ;
  assign n1140 = x3 & ~n1139 ;
  assign n1141 = n1136 & ~n1140 ;
  assign n1142 = x2 | n1141 ;
  assign n1143 = ( x4 & n68 ) | ( x4 & ~n764 ) | ( n68 & ~n764 ) ;
  assign n1144 = ~x3 & n1143 ;
  assign n1145 = x1 & n1144 ;
  assign n1146 = ( x1 & x7 ) | ( x1 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n1147 = ( x5 & ~x8 ) | ( x5 & n1146 ) | ( ~x8 & n1146 ) ;
  assign n1148 = x8 & n1147 ;
  assign n1149 = n1147 & ~n1148 ;
  assign n1150 = ( x8 & ~n1148 ) | ( x8 & n1149 ) | ( ~n1148 & n1149 ) ;
  assign n1151 = ( ~x3 & x4 ) | ( ~x3 & n1150 ) | ( x4 & n1150 ) ;
  assign n1152 = ( n60 & ~n1145 ) | ( n60 & n1151 ) | ( ~n1145 & n1151 ) ;
  assign n1153 = x0 | n1152 ;
  assign n1154 = x2 & n1153 ;
  assign n1155 = n1142 & ~n1154 ;
  assign n1156 = ( n38 & ~n596 ) | ( n38 & n729 ) | ( ~n596 & n729 ) ;
  assign n1157 = x3 & ~n192 ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1159 = ~x5 & n920 ;
  assign n1160 = ( ~n192 & n1157 ) | ( ~n192 & n1159 ) | ( n1157 & n1159 ) ;
  assign n1161 = ( x4 & n1158 ) | ( x4 & n1160 ) | ( n1158 & n1160 ) ;
  assign n1162 = x2 | n1161 ;
  assign n1163 = ~x5 & n729 ;
  assign n1164 = n26 & n1163 ;
  assign n1165 = x2 & ~n1164 ;
  assign n1166 = n1162 & ~n1165 ;
  assign n1167 = ( x6 & x7 ) | ( x6 & n83 ) | ( x7 & n83 ) ;
  assign n1168 = ( x6 & ~x8 ) | ( x6 & n83 ) | ( ~x8 & n83 ) ;
  assign n1169 = ( n20 & ~n1167 ) | ( n20 & n1168 ) | ( ~n1167 & n1168 ) ;
  assign n1170 = x5 & n1169 ;
  assign n1171 = x4 & n884 ;
  assign n1172 = x5 | n1171 ;
  assign n1173 = ~n1170 & n1172 ;
  assign n1174 = x2 & ~n1173 ;
  assign n1175 = n22 & n575 ;
  assign n1176 = x2 | n1175 ;
  assign n1177 = ~n1174 & n1176 ;
  assign n1178 = ( x2 & x4 ) | ( x2 & x7 ) | ( x4 & x7 ) ;
  assign n1179 = ( x2 & x3 ) | ( x2 & ~n1178 ) | ( x3 & ~n1178 ) ;
  assign n1180 = ( x4 & x7 ) | ( x4 & ~n1179 ) | ( x7 & ~n1179 ) ;
  assign n1181 = ~n1178 & n1180 ;
  assign n1182 = ( n1179 & n1180 ) | ( n1179 & n1181 ) | ( n1180 & n1181 ) ;
  assign n1183 = x5 & n49 ;
  assign n1184 = n1182 & n1183 ;
  assign n1185 = ( n1163 & n1182 ) | ( n1163 & n1184 ) | ( n1182 & n1184 ) ;
  assign n1186 = ( ~x3 & n1177 ) | ( ~x3 & n1185 ) | ( n1177 & n1185 ) ;
  assign n1187 = x2 & ~x6 ;
  assign n1188 = x7 & n53 ;
  assign n1189 = ( n572 & n1187 ) | ( n572 & ~n1188 ) | ( n1187 & ~n1188 ) ;
  assign n1190 = ( x2 & x4 ) | ( x2 & ~x6 ) | ( x4 & ~x6 ) ;
  assign n1191 = ( x2 & ~x7 ) | ( x2 & n1190 ) | ( ~x7 & n1190 ) ;
  assign n1192 = x2 & ~n1191 ;
  assign n1193 = n1191 | n1192 ;
  assign n1194 = ( ~x2 & n1192 ) | ( ~x2 & n1193 ) | ( n1192 & n1193 ) ;
  assign n1195 = x8 | n1194 ;
  assign n1196 = ( n1189 & n1194 ) | ( n1189 & n1195 ) | ( n1194 & n1195 ) ;
  assign n1197 = x5 | n1196 ;
  assign n1198 = ( x6 & x7 ) | ( x6 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n1199 = ( x2 & ~x6 ) | ( x2 & x8 ) | ( ~x6 & x8 ) ;
  assign n1200 = x7 & ~n1199 ;
  assign n1201 = n1198 & ~n1200 ;
  assign n1202 = ~x4 & n1201 ;
  assign n1203 = x5 & ~n1202 ;
  assign n1204 = n1197 & ~n1203 ;
  assign n1205 = ( x3 & n1185 ) | ( x3 & n1204 ) | ( n1185 & n1204 ) ;
  assign n1206 = n1186 | n1205 ;
  assign n1207 = x0 & n22 ;
  assign n1208 = ( n66 & ~n451 ) | ( n66 & n1207 ) | ( ~n451 & n1207 ) ;
  assign n1209 = ~n66 & n1208 ;
  assign n1210 = ( ~n1166 & n1206 ) | ( ~n1166 & n1209 ) | ( n1206 & n1209 ) ;
  assign n1211 = x0 & ~n1209 ;
  assign n1212 = ( n1166 & n1210 ) | ( n1166 & ~n1211 ) | ( n1210 & ~n1211 ) ;
  assign n1213 = x1 | n1212 ;
  assign n1214 = ( x2 & ~x4 ) | ( x2 & x5 ) | ( ~x4 & x5 ) ;
  assign n1215 = ( x2 & ~x7 ) | ( x2 & n1214 ) | ( ~x7 & n1214 ) ;
  assign n1216 = x2 & ~n1215 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = ( ~x2 & n1216 ) | ( ~x2 & n1217 ) | ( n1216 & n1217 ) ;
  assign n1219 = x8 & n1218 ;
  assign n1220 = ( x7 & n539 ) | ( x7 & ~n764 ) | ( n539 & ~n764 ) ;
  assign n1221 = ( x2 & ~x7 ) | ( x2 & n764 ) | ( ~x7 & n764 ) ;
  assign n1222 = ( ~x2 & n1220 ) | ( ~x2 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1223 = x8 | n1222 ;
  assign n1224 = ( ~x8 & n1219 ) | ( ~x8 & n1223 ) | ( n1219 & n1223 ) ;
  assign n1225 = x3 & ~n1224 ;
  assign n1226 = ( x4 & ~x5 ) | ( x4 & x8 ) | ( ~x5 & x8 ) ;
  assign n1227 = ~x2 & n1226 ;
  assign n1228 = ( n424 & n695 ) | ( n424 & ~n1227 ) | ( n695 & ~n1227 ) ;
  assign n1229 = x7 | n1228 ;
  assign n1230 = ~x3 & n1229 ;
  assign n1231 = n1225 | n1230 ;
  assign n1232 = x6 & ~n1231 ;
  assign n1233 = ( x2 & x5 ) | ( x2 & ~n488 ) | ( x5 & ~n488 ) ;
  assign n1234 = ( ~x5 & x7 ) | ( ~x5 & n1233 ) | ( x7 & n1233 ) ;
  assign n1235 = n488 | n1234 ;
  assign n1236 = ( ~x2 & n1233 ) | ( ~x2 & n1235 ) | ( n1233 & n1235 ) ;
  assign n1237 = x3 & n1236 ;
  assign n1238 = ( x5 & x7 ) | ( x5 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n1239 = x8 & n1238 ;
  assign n1240 = ( ~n738 & n1238 ) | ( ~n738 & n1239 ) | ( n1238 & n1239 ) ;
  assign n1241 = ~x2 & n1240 ;
  assign n1242 = x3 | n1241 ;
  assign n1243 = ~n1237 & n1242 ;
  assign n1244 = x4 | n1243 ;
  assign n1245 = ( x2 & x3 ) | ( x2 & ~n738 ) | ( x3 & ~n738 ) ;
  assign n1246 = ( ~x2 & x5 ) | ( ~x2 & n1245 ) | ( x5 & n1245 ) ;
  assign n1247 = ( ~x3 & x7 ) | ( ~x3 & n1246 ) | ( x7 & n1246 ) ;
  assign n1248 = n1245 & n1247 ;
  assign n1249 = ~x8 & n1248 ;
  assign n1250 = x4 & ~n1249 ;
  assign n1251 = n1244 & ~n1250 ;
  assign n1252 = x6 | n1251 ;
  assign n1253 = ( ~x6 & n1232 ) | ( ~x6 & n1252 ) | ( n1232 & n1252 ) ;
  assign n1254 = ~x0 & n1253 ;
  assign n1255 = x1 & ~n1254 ;
  assign n1256 = n1213 & ~n1255 ;
  assign n1257 = n1155 | n1256 ;
  assign n1258 = ( ~n1122 & n1123 ) | ( ~n1122 & n1257 ) | ( n1123 & n1257 ) ;
  assign n1259 = ~x0 & x2 ;
  assign n1260 = x0 & ~x5 ;
  assign n1261 = ( ~n155 & n1259 ) | ( ~n155 & n1260 ) | ( n1259 & n1260 ) ;
  assign n1262 = x6 | n1261 ;
  assign n1263 = ~x0 & x4 ;
  assign n1264 = ( n285 & n1259 ) | ( n285 & ~n1263 ) | ( n1259 & ~n1263 ) ;
  assign n1265 = ~x5 & n1264 ;
  assign n1266 = x6 & ~n1265 ;
  assign n1267 = n1262 & ~n1266 ;
  assign n1268 = x1 | n1267 ;
  assign n1269 = x6 & ~n539 ;
  assign n1270 = ( n52 & n118 ) | ( n52 & ~n1269 ) | ( n118 & ~n1269 ) ;
  assign n1271 = ~x0 & n1270 ;
  assign n1272 = x1 & ~n1271 ;
  assign n1273 = n1268 & ~n1272 ;
  assign n1274 = x3 | n1273 ;
  assign n1275 = ( x1 & x4 ) | ( x1 & ~n764 ) | ( x4 & ~n764 ) ;
  assign n1276 = ( x1 & x2 ) | ( x1 & ~n764 ) | ( x2 & ~n764 ) ;
  assign n1277 = ( n539 & n1275 ) | ( n539 & ~n1276 ) | ( n1275 & ~n1276 ) ;
  assign n1278 = ~x6 & n22 ;
  assign n1279 = n511 & n1278 ;
  assign n1280 = x6 | n1279 ;
  assign n1281 = ( n1277 & n1279 ) | ( n1277 & n1280 ) | ( n1279 & n1280 ) ;
  assign n1282 = ~x0 & n1281 ;
  assign n1283 = x3 & ~n1282 ;
  assign n1284 = n1274 & ~n1283 ;
  assign n1285 = n1258 | n1284 ;
  assign n1286 = ( n21 & n1258 ) | ( n21 & n1285 ) | ( n1258 & n1285 ) ;
  assign n1287 = x2 | x6 ;
  assign n1288 = ( ~n201 & n330 ) | ( ~n201 & n1287 ) | ( n330 & n1287 ) ;
  assign n1289 = x1 & ~n1288 ;
  assign n1290 = ~x0 & n1289 ;
  assign n1291 = ( x2 & n98 ) | ( x2 & n463 ) | ( n98 & n463 ) ;
  assign n1292 = ~x2 & n1291 ;
  assign n1293 = x4 & ~n15 ;
  assign n1294 = ( x6 & x7 ) | ( x6 & n1293 ) | ( x7 & n1293 ) ;
  assign n1295 = ~x7 & n1294 ;
  assign n1296 = n105 | n1295 ;
  assign n1297 = ( n1101 & n1295 ) | ( n1101 & n1296 ) | ( n1295 & n1296 ) ;
  assign n1298 = x0 & n1297 ;
  assign n1299 = ~x4 & n320 ;
  assign n1300 = ~n566 & n1299 ;
  assign n1301 = ( x6 & ~x7 ) | ( x6 & n1083 ) | ( ~x7 & n1083 ) ;
  assign n1302 = ( x2 & x6 ) | ( x2 & ~n1083 ) | ( x6 & ~n1083 ) ;
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = ( x0 & x8 ) | ( x0 & n1303 ) | ( x8 & n1303 ) ;
  assign n1305 = x0 & x4 ;
  assign n1306 = ( x2 & ~n566 ) | ( x2 & n1305 ) | ( ~n566 & n1305 ) ;
  assign n1307 = ~x2 & n1306 ;
  assign n1308 = x8 & n1307 ;
  assign n1309 = ( ~x0 & n1304 ) | ( ~x0 & n1308 ) | ( n1304 & n1308 ) ;
  assign n1310 = ( ~x4 & x6 ) | ( ~x4 & x7 ) | ( x6 & x7 ) ;
  assign n1311 = ( ~x4 & x6 ) | ( ~x4 & x8 ) | ( x6 & x8 ) ;
  assign n1312 = n1310 & ~n1311 ;
  assign n1313 = ( ~x0 & n1309 ) | ( ~x0 & n1312 ) | ( n1309 & n1312 ) ;
  assign n1314 = x2 & ~n1313 ;
  assign n1315 = ( x2 & n1309 ) | ( x2 & ~n1314 ) | ( n1309 & ~n1314 ) ;
  assign n1316 = x1 | n1315 ;
  assign n1317 = ( ~x2 & x8 ) | ( ~x2 & n446 ) | ( x8 & n446 ) ;
  assign n1318 = n487 & n1317 ;
  assign n1319 = ~x0 & n1318 ;
  assign n1320 = x1 & ~n1319 ;
  assign n1321 = n1316 & ~n1320 ;
  assign n1322 = n1300 | n1321 ;
  assign n1323 = ( n1297 & ~n1298 ) | ( n1297 & n1322 ) | ( ~n1298 & n1322 ) ;
  assign n1324 = ( ~n1290 & n1292 ) | ( ~n1290 & n1323 ) | ( n1292 & n1323 ) ;
  assign n1325 = n21 & ~n1323 ;
  assign n1326 = ( n1290 & n1324 ) | ( n1290 & ~n1325 ) | ( n1324 & ~n1325 ) ;
  assign n1327 = x3 & n1326 ;
  assign n1328 = ( x1 & x2 ) | ( x1 & x4 ) | ( x2 & x4 ) ;
  assign n1329 = ( x2 & x6 ) | ( x2 & ~n1328 ) | ( x6 & ~n1328 ) ;
  assign n1330 = ( x1 & x4 ) | ( x1 & ~n1329 ) | ( x4 & ~n1329 ) ;
  assign n1331 = n1328 & ~n1330 ;
  assign n1332 = ( n1329 & n1330 ) | ( n1329 & ~n1331 ) | ( n1330 & ~n1331 ) ;
  assign n1333 = ( ~x7 & x8 ) | ( ~x7 & n1332 ) | ( x8 & n1332 ) ;
  assign n1334 = ~x2 & x6 ;
  assign n1335 = ( x2 & x4 ) | ( x2 & n1334 ) | ( x4 & n1334 ) ;
  assign n1336 = ( x1 & x4 ) | ( x1 & n1334 ) | ( x4 & n1334 ) ;
  assign n1337 = ( n511 & n1335 ) | ( n511 & ~n1336 ) | ( n1335 & ~n1336 ) ;
  assign n1338 = ( x7 & x8 ) | ( x7 & ~n1337 ) | ( x8 & ~n1337 ) ;
  assign n1339 = n1333 | n1338 ;
  assign n1340 = ( ~x2 & x4 ) | ( ~x2 & n908 ) | ( x4 & n908 ) ;
  assign n1341 = ( x4 & x6 ) | ( x4 & ~n908 ) | ( x6 & ~n908 ) ;
  assign n1342 = n1340 & ~n1341 ;
  assign n1343 = ( x1 & x8 ) | ( x1 & ~n1342 ) | ( x8 & ~n1342 ) ;
  assign n1344 = ( x2 & x4 ) | ( x2 & ~n72 ) | ( x4 & ~n72 ) ;
  assign n1345 = ( ~x1 & x4 ) | ( ~x1 & n72 ) | ( x4 & n72 ) ;
  assign n1346 = n1344 & ~n1345 ;
  assign n1347 = x8 & n1346 ;
  assign n1348 = ( n1342 & n1343 ) | ( n1342 & n1347 ) | ( n1343 & n1347 ) ;
  assign n1349 = n1339 & n1348 ;
  assign n1350 = ~x0 & x3 ;
  assign n1351 = ( ~n1339 & n1349 ) | ( ~n1339 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1352 = ( ~x1 & n26 ) | ( ~x1 & n587 ) | ( n26 & n587 ) ;
  assign n1353 = x1 & n936 ;
  assign n1354 = ( n26 & ~n1352 ) | ( n26 & n1353 ) | ( ~n1352 & n1353 ) ;
  assign n1355 = ( x0 & ~x2 ) | ( x0 & n1354 ) | ( ~x2 & n1354 ) ;
  assign n1356 = x1 | x3 ;
  assign n1357 = x0 & ~n1356 ;
  assign n1358 = x4 & n596 ;
  assign n1359 = n1357 & n1358 ;
  assign n1360 = ~x2 & n1359 ;
  assign n1361 = ( ~x0 & n1355 ) | ( ~x0 & n1360 ) | ( n1355 & n1360 ) ;
  assign n1362 = ( n106 & n192 ) | ( n106 & n1361 ) | ( n192 & n1361 ) ;
  assign n1363 = n596 & ~n1362 ;
  assign n1364 = ( n596 & n1361 ) | ( n596 & ~n1363 ) | ( n1361 & ~n1363 ) ;
  assign n1365 = n21 & n1364 ;
  assign n1366 = n99 & ~n451 ;
  assign n1367 = n118 & n1366 ;
  assign n1368 = ~x4 & n596 ;
  assign n1369 = ( x1 & n227 ) | ( x1 & n1368 ) | ( n227 & n1368 ) ;
  assign n1370 = ~x1 & n1369 ;
  assign n1371 = ( x1 & ~x3 ) | ( x1 & x4 ) | ( ~x3 & x4 ) ;
  assign n1372 = ( x1 & x6 ) | ( x1 & ~n1371 ) | ( x6 & ~n1371 ) ;
  assign n1373 = ( x3 & ~x4 ) | ( x3 & n1372 ) | ( ~x4 & n1372 ) ;
  assign n1374 = n1371 | n1373 ;
  assign n1375 = ( ~n1372 & n1373 ) | ( ~n1372 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1376 = ( x2 & ~n1370 ) | ( x2 & n1375 ) | ( ~n1370 & n1375 ) ;
  assign n1377 = ~x5 & n1376 ;
  assign n1378 = ( x5 & ~n1370 ) | ( x5 & n1377 ) | ( ~n1370 & n1377 ) ;
  assign n1379 = ( x0 & ~n1367 ) | ( x0 & n1378 ) | ( ~n1367 & n1378 ) ;
  assign n1380 = x8 & n1379 ;
  assign n1381 = ( x8 & n1367 ) | ( x8 & ~n1380 ) | ( n1367 & ~n1380 ) ;
  assign n1382 = x1 & ~n511 ;
  assign n1383 = n452 & n1382 ;
  assign n1384 = ~x4 & n920 ;
  assign n1385 = ( ~n511 & n1382 ) | ( ~n511 & n1384 ) | ( n1382 & n1384 ) ;
  assign n1386 = ( ~x2 & n1383 ) | ( ~x2 & n1385 ) | ( n1383 & n1385 ) ;
  assign n1387 = ( ~x3 & n376 ) | ( ~x3 & n672 ) | ( n376 & n672 ) ;
  assign n1388 = n1386 & n1387 ;
  assign n1389 = ( x2 & x3 ) | ( x2 & x5 ) | ( x3 & x5 ) ;
  assign n1390 = ( x3 & ~x4 ) | ( x3 & n1389 ) | ( ~x4 & n1389 ) ;
  assign n1391 = x3 & ~n1390 ;
  assign n1392 = n1390 | n1391 ;
  assign n1393 = ( ~x3 & n1391 ) | ( ~x3 & n1392 ) | ( n1391 & n1392 ) ;
  assign n1394 = ( x1 & ~x8 ) | ( x1 & n1393 ) | ( ~x8 & n1393 ) ;
  assign n1395 = x8 & n1394 ;
  assign n1396 = ( x1 & x6 ) | ( x1 & ~n1395 ) | ( x6 & ~n1395 ) ;
  assign n1397 = ( n1394 & n1395 ) | ( n1394 & ~n1396 ) | ( n1395 & ~n1396 ) ;
  assign n1398 = ( x2 & x3 ) | ( x2 & ~x4 ) | ( x3 & ~x4 ) ;
  assign n1399 = ( x4 & x6 ) | ( x4 & n1398 ) | ( x6 & n1398 ) ;
  assign n1400 = ( x2 & x3 ) | ( x2 & n1399 ) | ( x3 & n1399 ) ;
  assign n1401 = ~n1398 & n1400 ;
  assign n1402 = ( ~n1399 & n1400 ) | ( ~n1399 & n1401 ) | ( n1400 & n1401 ) ;
  assign n1403 = x5 & ~n1402 ;
  assign n1404 = ~x3 & n446 ;
  assign n1405 = x5 | n1404 ;
  assign n1406 = ~n1403 & n1405 ;
  assign n1407 = x1 | n1406 ;
  assign n1408 = ~n66 & n1358 ;
  assign n1409 = x1 & ~n1408 ;
  assign n1410 = n1407 & ~n1409 ;
  assign n1411 = ~x8 & n1410 ;
  assign n1412 = ( x2 & x6 ) | ( x2 & n111 ) | ( x6 & n111 ) ;
  assign n1413 = ( x5 & x6 ) | ( x5 & ~n1412 ) | ( x6 & ~n1412 ) ;
  assign n1414 = n111 | n1413 ;
  assign n1415 = ( x2 & ~n1412 ) | ( x2 & n1414 ) | ( ~n1412 & n1414 ) ;
  assign n1416 = ( ~x1 & x3 ) | ( ~x1 & n1415 ) | ( x3 & n1415 ) ;
  assign n1417 = n430 & ~n587 ;
  assign n1418 = ~x1 & n1417 ;
  assign n1419 = ( ~n1415 & n1416 ) | ( ~n1415 & n1418 ) | ( n1416 & n1418 ) ;
  assign n1420 = x3 & x6 ;
  assign n1421 = ( ~x2 & x5 ) | ( ~x2 & n1420 ) | ( x5 & n1420 ) ;
  assign n1422 = ( x5 & x6 ) | ( x5 & ~n1420 ) | ( x6 & ~n1420 ) ;
  assign n1423 = ( ~x2 & x3 ) | ( ~x2 & n1422 ) | ( x3 & n1422 ) ;
  assign n1424 = ~n1421 & n1423 ;
  assign n1425 = ( ~x1 & x4 ) | ( ~x1 & n1424 ) | ( x4 & n1424 ) ;
  assign n1426 = ( ~x5 & n587 ) | ( ~x5 & n825 ) | ( n587 & n825 ) ;
  assign n1427 = ( x2 & n26 ) | ( x2 & n1426 ) | ( n26 & n1426 ) ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = x1 & n1428 ;
  assign n1430 = ( n1424 & ~n1425 ) | ( n1424 & n1429 ) | ( ~n1425 & n1429 ) ;
  assign n1431 = n1419 | n1430 ;
  assign n1432 = x8 & n1431 ;
  assign n1433 = n1411 | n1432 ;
  assign n1434 = n1397 | n1433 ;
  assign n1435 = ( n1386 & ~n1388 ) | ( n1386 & n1434 ) | ( ~n1388 & n1434 ) ;
  assign n1436 = ( ~x0 & x7 ) | ( ~x0 & n1435 ) | ( x7 & n1435 ) ;
  assign n1437 = ( x1 & x3 ) | ( x1 & x6 ) | ( x3 & x6 ) ;
  assign n1438 = ( x3 & n596 ) | ( x3 & ~n1437 ) | ( n596 & ~n1437 ) ;
  assign n1439 = ( ~x5 & n1437 ) | ( ~x5 & n1438 ) | ( n1437 & n1438 ) ;
  assign n1440 = ( ~x3 & n1438 ) | ( ~x3 & n1439 ) | ( n1438 & n1439 ) ;
  assign n1441 = ( ~x2 & x8 ) | ( ~x2 & n1440 ) | ( x8 & n1440 ) ;
  assign n1442 = x6 | n15 ;
  assign n1443 = ( x3 & x5 ) | ( x3 & ~n1442 ) | ( x5 & ~n1442 ) ;
  assign n1444 = ~x3 & n1443 ;
  assign n1445 = ~x8 & n1444 ;
  assign n1446 = ( n1440 & ~n1441 ) | ( n1440 & n1445 ) | ( ~n1441 & n1445 ) ;
  assign n1447 = ( ~x1 & n1183 ) | ( ~x1 & n1446 ) | ( n1183 & n1446 ) ;
  assign n1448 = n842 & ~n1447 ;
  assign n1449 = ( n842 & n1446 ) | ( n842 & ~n1448 ) | ( n1446 & ~n1448 ) ;
  assign n1450 = ( x3 & x8 ) | ( x3 & ~n879 ) | ( x8 & ~n879 ) ;
  assign n1451 = ( x3 & x5 ) | ( x3 & ~n879 ) | ( x5 & ~n879 ) ;
  assign n1452 = ( n613 & n1450 ) | ( n613 & ~n1451 ) | ( n1450 & ~n1451 ) ;
  assign n1453 = ( x2 & x6 ) | ( x2 & n1452 ) | ( x6 & n1452 ) ;
  assign n1454 = ( x1 & ~x2 ) | ( x1 & n1453 ) | ( ~x2 & n1453 ) ;
  assign n1455 = ( x1 & x6 ) | ( x1 & ~n1453 ) | ( x6 & ~n1453 ) ;
  assign n1456 = n1454 & ~n1455 ;
  assign n1457 = ( ~x4 & n1449 ) | ( ~x4 & n1456 ) | ( n1449 & n1456 ) ;
  assign n1458 = ( x3 & ~x6 ) | ( x3 & n1287 ) | ( ~x6 & n1287 ) ;
  assign n1459 = ( x3 & ~x5 ) | ( x3 & n1287 ) | ( ~x5 & n1287 ) ;
  assign n1460 = ( n825 & ~n1458 ) | ( n825 & n1459 ) | ( ~n1458 & n1459 ) ;
  assign n1461 = x1 & x8 ;
  assign n1462 = x8 & ~n1461 ;
  assign n1463 = n1460 & n1462 ;
  assign n1464 = ( x2 & x5 ) | ( x2 & x6 ) | ( x5 & x6 ) ;
  assign n1465 = ~x3 & x6 ;
  assign n1466 = ( n1389 & ~n1464 ) | ( n1389 & n1465 ) | ( ~n1464 & n1465 ) ;
  assign n1467 = ( ~n1461 & n1462 ) | ( ~n1461 & n1466 ) | ( n1462 & n1466 ) ;
  assign n1468 = ( x1 & n1463 ) | ( x1 & n1467 ) | ( n1463 & n1467 ) ;
  assign n1469 = ( x4 & n1456 ) | ( x4 & n1468 ) | ( n1456 & n1468 ) ;
  assign n1470 = n1457 | n1469 ;
  assign n1471 = ( x0 & x7 ) | ( x0 & ~n1470 ) | ( x7 & ~n1470 ) ;
  assign n1472 = n1436 & ~n1471 ;
  assign n1473 = ( n99 & n258 ) | ( n99 & n1472 ) | ( n258 & n1472 ) ;
  assign n1474 = n67 & ~n1473 ;
  assign n1475 = ( n67 & n1472 ) | ( n67 & ~n1474 ) | ( n1472 & ~n1474 ) ;
  assign n1476 = n1381 | n1475 ;
  assign n1477 = ( n1364 & ~n1365 ) | ( n1364 & n1476 ) | ( ~n1365 & n1476 ) ;
  assign n1478 = n1351 | n1477 ;
  assign n1479 = ( n1326 & ~n1327 ) | ( n1326 & n1478 ) | ( ~n1327 & n1478 ) ;
  assign n1480 = ~x3 & n347 ;
  assign n1481 = ( x1 & ~x4 ) | ( x1 & n1480 ) | ( ~x4 & n1480 ) ;
  assign n1482 = ( n347 & n1480 ) | ( n347 & n1481 ) | ( n1480 & n1481 ) ;
  assign n1483 = x6 & n1482 ;
  assign n1484 = x1 | x8 ;
  assign n1485 = ( n689 & ~n911 ) | ( n689 & n1484 ) | ( ~n911 & n1484 ) ;
  assign n1486 = ( x3 & x6 ) | ( x3 & ~n1485 ) | ( x6 & ~n1485 ) ;
  assign n1487 = ( ~n1420 & n1483 ) | ( ~n1420 & n1486 ) | ( n1483 & n1486 ) ;
  assign n1488 = x5 & ~n1487 ;
  assign n1489 = ( x4 & x6 ) | ( x4 & ~x8 ) | ( x6 & ~x8 ) ;
  assign n1490 = ~x4 & n1489 ;
  assign n1491 = ( ~x3 & x8 ) | ( ~x3 & n1490 ) | ( x8 & n1490 ) ;
  assign n1492 = ( n1489 & n1490 ) | ( n1489 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1493 = x1 & n1492 ;
  assign n1494 = x5 | n1493 ;
  assign n1495 = ~n1488 & n1494 ;
  assign n1496 = ( x2 & ~x7 ) | ( x2 & n1495 ) | ( ~x7 & n1495 ) ;
  assign n1497 = x3 & ~n38 ;
  assign n1498 = ( x5 & x6 ) | ( x5 & ~n38 ) | ( x6 & ~n38 ) ;
  assign n1499 = ( x3 & n587 ) | ( x3 & ~n1498 ) | ( n587 & ~n1498 ) ;
  assign n1500 = ( ~x3 & n1497 ) | ( ~x3 & n1499 ) | ( n1497 & n1499 ) ;
  assign n1501 = x1 | n1500 ;
  assign n1502 = x5 & ~n451 ;
  assign n1503 = ~x3 & n1502 ;
  assign n1504 = x1 & ~n1503 ;
  assign n1505 = n1501 & ~n1504 ;
  assign n1506 = x4 & n1505 ;
  assign n1507 = ( x1 & ~x3 ) | ( x1 & x6 ) | ( ~x3 & x6 ) ;
  assign n1508 = ( x3 & x5 ) | ( x3 & n1507 ) | ( x5 & n1507 ) ;
  assign n1509 = x3 & n1507 ;
  assign n1510 = x5 | n1507 ;
  assign n1511 = ( ~n1508 & n1509 ) | ( ~n1508 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = x8 & ~n1511 ;
  assign n1513 = ( n37 & n74 ) | ( n37 & ~n576 ) | ( n74 & ~n576 ) ;
  assign n1514 = x6 & n1513 ;
  assign n1515 = x8 | n1514 ;
  assign n1516 = ~n1512 & n1515 ;
  assign n1517 = x4 | n1516 ;
  assign n1518 = ( ~x4 & n1506 ) | ( ~x4 & n1517 ) | ( n1506 & n1517 ) ;
  assign n1519 = ( x2 & x7 ) | ( x2 & n1518 ) | ( x7 & n1518 ) ;
  assign n1520 = n1496 & n1519 ;
  assign n1521 = x0 & n1520 ;
  assign n1522 = n1116 & ~n1356 ;
  assign n1523 = ( x3 & n566 ) | ( x3 & n911 ) | ( n566 & n911 ) ;
  assign n1524 = ~n566 & n1523 ;
  assign n1525 = n1522 | n1524 ;
  assign n1526 = ( ~x0 & n1522 ) | ( ~x0 & n1525 ) | ( n1522 & n1525 ) ;
  assign n1527 = ( x2 & n614 ) | ( x2 & n1526 ) | ( n614 & n1526 ) ;
  assign n1528 = ( n37 & ~n306 ) | ( n37 & n695 ) | ( ~n306 & n695 ) ;
  assign n1529 = x7 & n1528 ;
  assign n1530 = x3 & x8 ;
  assign n1531 = ( x4 & ~x5 ) | ( x4 & n1530 ) | ( ~x5 & n1530 ) ;
  assign n1532 = ( ~x3 & x5 ) | ( ~x3 & n1531 ) | ( x5 & n1531 ) ;
  assign n1533 = ( x4 & x8 ) | ( x4 & ~n1532 ) | ( x8 & ~n1532 ) ;
  assign n1534 = ~n1531 & n1533 ;
  assign n1535 = x7 | n1534 ;
  assign n1536 = x5 & n187 ;
  assign n1537 = x5 | n879 ;
  assign n1538 = ~n1536 & n1537 ;
  assign n1539 = x3 & ~n1538 ;
  assign n1540 = x7 & ~n1539 ;
  assign n1541 = n1535 & ~n1540 ;
  assign n1542 = ~x3 & n176 ;
  assign n1543 = x0 & n1542 ;
  assign n1544 = ( ~n1529 & n1541 ) | ( ~n1529 & n1543 ) | ( n1541 & n1543 ) ;
  assign n1545 = x0 & ~n1543 ;
  assign n1546 = ( n1529 & n1544 ) | ( n1529 & ~n1545 ) | ( n1544 & ~n1545 ) ;
  assign n1547 = x6 & ~n1546 ;
  assign n1548 = ( x3 & ~n785 ) | ( x3 & n879 ) | ( ~n785 & n879 ) ;
  assign n1549 = ( ~x3 & x7 ) | ( ~x3 & n1548 ) | ( x7 & n1548 ) ;
  assign n1550 = ( ~x4 & n879 ) | ( ~x4 & n1549 ) | ( n879 & n1549 ) ;
  assign n1551 = ( ~n879 & n1548 ) | ( ~n879 & n1550 ) | ( n1548 & n1550 ) ;
  assign n1552 = x5 & n1551 ;
  assign n1553 = ( x3 & x7 ) | ( x3 & x8 ) | ( x7 & x8 ) ;
  assign n1554 = ~x3 & n1553 ;
  assign n1555 = ( ~n68 & n1553 ) | ( ~n68 & n1554 ) | ( n1553 & n1554 ) ;
  assign n1556 = x4 & n1555 ;
  assign n1557 = x5 | n1556 ;
  assign n1558 = ~n1552 & n1557 ;
  assign n1559 = ~x0 & n1558 ;
  assign n1560 = x6 | n1559 ;
  assign n1561 = ~n1547 & n1560 ;
  assign n1562 = x1 | n1561 ;
  assign n1563 = ( x3 & ~x4 ) | ( x3 & x7 ) | ( ~x4 & x7 ) ;
  assign n1564 = ( x3 & ~x6 ) | ( x3 & n1563 ) | ( ~x6 & n1563 ) ;
  assign n1565 = x3 & ~n1564 ;
  assign n1566 = n1564 | n1565 ;
  assign n1567 = ( ~x3 & n1565 ) | ( ~x3 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1568 = x8 & n1567 ;
  assign n1569 = ( x4 & x6 ) | ( x4 & ~x7 ) | ( x6 & ~x7 ) ;
  assign n1570 = x4 & ~n1569 ;
  assign n1571 = ( n551 & n1569 ) | ( n551 & ~n1570 ) | ( n1569 & ~n1570 ) ;
  assign n1572 = ~x8 & n1571 ;
  assign n1573 = ( x8 & ~n1568 ) | ( x8 & n1572 ) | ( ~n1568 & n1572 ) ;
  assign n1574 = x5 & ~n1573 ;
  assign n1575 = x3 | x7 ;
  assign n1576 = x6 & n1575 ;
  assign n1577 = ( n68 & n729 ) | ( n68 & ~n1576 ) | ( n729 & ~n1576 ) ;
  assign n1578 = ~x4 & n1577 ;
  assign n1579 = ( n10 & n451 ) | ( n10 & ~n572 ) | ( n451 & ~n572 ) ;
  assign n1580 = ( x3 & x4 ) | ( x3 & n1579 ) | ( x4 & n1579 ) ;
  assign n1581 = ( n95 & n1578 ) | ( n95 & ~n1580 ) | ( n1578 & ~n1580 ) ;
  assign n1582 = x5 | n1581 ;
  assign n1583 = ( ~x5 & n1574 ) | ( ~x5 & n1582 ) | ( n1574 & n1582 ) ;
  assign n1584 = ~x0 & n1583 ;
  assign n1585 = x1 & ~n1584 ;
  assign n1586 = n1562 & ~n1585 ;
  assign n1587 = ~x2 & n1586 ;
  assign n1588 = ( n1526 & ~n1527 ) | ( n1526 & n1587 ) | ( ~n1527 & n1587 ) ;
  assign n1589 = ~n384 & n1190 ;
  assign n1590 = ( ~x0 & x1 ) | ( ~x0 & n1589 ) | ( x1 & n1589 ) ;
  assign n1591 = x4 & n52 ;
  assign n1592 = n511 & n1591 ;
  assign n1593 = ~x0 & n1592 ;
  assign n1594 = ( ~x1 & n1590 ) | ( ~x1 & n1593 ) | ( n1590 & n1593 ) ;
  assign n1595 = ( ~n106 & n320 ) | ( ~n106 & n1594 ) | ( n320 & n1594 ) ;
  assign n1596 = ( n22 & n52 ) | ( n22 & ~n463 ) | ( n52 & ~n463 ) ;
  assign n1597 = n1594 | n1596 ;
  assign n1598 = ( n106 & n1595 ) | ( n106 & n1597 ) | ( n1595 & n1597 ) ;
  assign n1599 = x8 | n1598 ;
  assign n1600 = ( x2 & ~x4 ) | ( x2 & x6 ) | ( ~x4 & x6 ) ;
  assign n1601 = ( x2 & ~x5 ) | ( x2 & n1600 ) | ( ~x5 & n1600 ) ;
  assign n1602 = x2 & ~n1601 ;
  assign n1603 = n1601 | n1602 ;
  assign n1604 = ( ~x2 & n1602 ) | ( ~x2 & n1603 ) | ( n1602 & n1603 ) ;
  assign n1605 = x1 & n1604 ;
  assign n1606 = ( x2 & ~x4 ) | ( x2 & n705 ) | ( ~x4 & n705 ) ;
  assign n1607 = ( x5 & x6 ) | ( x5 & n1606 ) | ( x6 & n1606 ) ;
  assign n1608 = n705 & ~n1607 ;
  assign n1609 = ( n1606 & ~n1607 ) | ( n1606 & n1608 ) | ( ~n1607 & n1608 ) ;
  assign n1610 = x1 | n1609 ;
  assign n1611 = ( ~x1 & n1605 ) | ( ~x1 & n1610 ) | ( n1605 & n1610 ) ;
  assign n1612 = ~x0 & n1611 ;
  assign n1613 = x8 & ~n1612 ;
  assign n1614 = n1599 & ~n1613 ;
  assign n1615 = x3 | n1614 ;
  assign n1616 = ( x2 & n911 ) | ( x2 & n1163 ) | ( n911 & n1163 ) ;
  assign n1617 = ~x2 & n1616 ;
  assign n1618 = ( x1 & x4 ) | ( x1 & x8 ) | ( x4 & x8 ) ;
  assign n1619 = ( x6 & x8 ) | ( x6 & n911 ) | ( x8 & n911 ) ;
  assign n1620 = n1618 & ~n1619 ;
  assign n1621 = ( x2 & n1617 ) | ( x2 & n1620 ) | ( n1617 & n1620 ) ;
  assign n1622 = x5 & ~n1621 ;
  assign n1623 = ( x5 & n1617 ) | ( x5 & ~n1622 ) | ( n1617 & ~n1622 ) ;
  assign n1624 = ~x0 & n1623 ;
  assign n1625 = x3 & ~n1624 ;
  assign n1626 = n1615 & ~n1625 ;
  assign n1627 = n1588 | n1626 ;
  assign n1628 = ( n1520 & ~n1521 ) | ( n1520 & n1627 ) | ( ~n1521 & n1627 ) ;
  assign n1629 = ( x1 & x3 ) | ( x1 & x7 ) | ( x3 & x7 ) ;
  assign n1630 = ( x1 & x4 ) | ( x1 & x7 ) | ( x4 & x7 ) ;
  assign n1631 = ( n60 & ~n1629 ) | ( n60 & n1630 ) | ( ~n1629 & n1630 ) ;
  assign n1632 = ( x2 & x8 ) | ( x2 & ~n1631 ) | ( x8 & ~n1631 ) ;
  assign n1633 = x1 & x3 ;
  assign n1634 = ( x4 & x8 ) | ( x4 & n1633 ) | ( x8 & n1633 ) ;
  assign n1635 = ~x8 & n1634 ;
  assign n1636 = x2 & n1635 ;
  assign n1637 = ( n1631 & n1632 ) | ( n1631 & n1636 ) | ( n1632 & n1636 ) ;
  assign n1638 = ( ~x3 & x4 ) | ( ~x3 & x8 ) | ( x4 & x8 ) ;
  assign n1639 = ( x3 & x7 ) | ( x3 & n1638 ) | ( x7 & n1638 ) ;
  assign n1640 = ( x4 & x8 ) | ( x4 & n1639 ) | ( x8 & n1639 ) ;
  assign n1641 = n1638 & ~n1640 ;
  assign n1642 = ( n1639 & ~n1640 ) | ( n1639 & n1641 ) | ( ~n1640 & n1641 ) ;
  assign n1643 = ( x1 & ~x2 ) | ( x1 & n1642 ) | ( ~x2 & n1642 ) ;
  assign n1644 = ( x3 & x4 ) | ( x3 & x8 ) | ( x4 & x8 ) ;
  assign n1645 = ( x4 & ~x7 ) | ( x4 & n1644 ) | ( ~x7 & n1644 ) ;
  assign n1646 = x4 & ~n1645 ;
  assign n1647 = n1645 | n1646 ;
  assign n1648 = ( ~x4 & n1646 ) | ( ~x4 & n1647 ) | ( n1646 & n1647 ) ;
  assign n1649 = ( x1 & x2 ) | ( x1 & ~n1648 ) | ( x2 & ~n1648 ) ;
  assign n1650 = n1643 & ~n1649 ;
  assign n1651 = ( x3 & ~x7 ) | ( x3 & n105 ) | ( ~x7 & n105 ) ;
  assign n1652 = ( x1 & x3 ) | ( x1 & ~n105 ) | ( x3 & ~n105 ) ;
  assign n1653 = ( x2 & ~x7 ) | ( x2 & n1652 ) | ( ~x7 & n1652 ) ;
  assign n1654 = ~n1651 & n1653 ;
  assign n1655 = ( x0 & n880 ) | ( x0 & n1654 ) | ( n880 & n1654 ) ;
  assign n1656 = ~x3 & x7 ;
  assign n1657 = ( x2 & n98 ) | ( x2 & n1656 ) | ( n98 & n1656 ) ;
  assign n1658 = ~x2 & n1657 ;
  assign n1659 = ~n880 & n1658 ;
  assign n1660 = ( n1654 & ~n1655 ) | ( n1654 & n1659 ) | ( ~n1655 & n1659 ) ;
  assign n1661 = ( ~n1637 & n1650 ) | ( ~n1637 & n1660 ) | ( n1650 & n1660 ) ;
  assign n1662 = x0 & ~n1660 ;
  assign n1663 = ( n1637 & n1661 ) | ( n1637 & ~n1662 ) | ( n1661 & ~n1662 ) ;
  assign n1664 = n1628 | n1663 ;
  assign n1665 = ( ~n1426 & n1628 ) | ( ~n1426 & n1664 ) | ( n1628 & n1664 ) ;
  assign n1666 = ( n95 & ~n118 ) | ( n95 & n786 ) | ( ~n118 & n786 ) ;
  assign n1667 = ( ~x3 & n95 ) | ( ~x3 & n1666 ) | ( n95 & n1666 ) ;
  assign n1668 = x1 & ~n1667 ;
  assign n1669 = ~x0 & n1668 ;
  assign n1670 = n377 & ~n1669 ;
  assign n1671 = ( n320 & n1669 ) | ( n320 & ~n1670 ) | ( n1669 & ~n1670 ) ;
  assign n1672 = n320 & n596 ;
  assign n1673 = n26 & n1672 ;
  assign n1674 = x5 | n57 ;
  assign n1675 = ( ~n764 & n911 ) | ( ~n764 & n1674 ) | ( n911 & n1674 ) ;
  assign n1676 = ( n22 & n330 ) | ( n22 & ~n825 ) | ( n330 & ~n825 ) ;
  assign n1677 = ( x1 & ~x2 ) | ( x1 & n1676 ) | ( ~x2 & n1676 ) ;
  assign n1678 = ~x1 & n1677 ;
  assign n1679 = ( x2 & n1677 ) | ( x2 & n1678 ) | ( n1677 & n1678 ) ;
  assign n1680 = x6 | n1679 ;
  assign n1681 = ( n1675 & n1679 ) | ( n1675 & n1680 ) | ( n1679 & n1680 ) ;
  assign n1682 = ( ~x0 & x3 ) | ( ~x0 & n1681 ) | ( x3 & n1681 ) ;
  assign n1683 = ( x1 & x4 ) | ( x1 & ~n15 ) | ( x4 & ~n15 ) ;
  assign n1684 = ( x4 & x5 ) | ( x4 & ~n15 ) | ( x5 & ~n15 ) ;
  assign n1685 = ( n576 & n1683 ) | ( n576 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1686 = ~x6 & n1685 ;
  assign n1687 = ( x1 & ~x2 ) | ( x1 & x6 ) | ( ~x2 & x6 ) ;
  assign n1688 = n1054 & n1687 ;
  assign n1689 = n1686 | n1688 ;
  assign n1690 = ( ~x4 & n1686 ) | ( ~x4 & n1689 ) | ( n1686 & n1689 ) ;
  assign n1691 = ( x0 & x3 ) | ( x0 & ~n1690 ) | ( x3 & ~n1690 ) ;
  assign n1692 = n1682 & ~n1691 ;
  assign n1693 = ( ~n21 & n1673 ) | ( ~n21 & n1692 ) | ( n1673 & n1692 ) ;
  assign n1694 = ~n1671 & n1693 ;
  assign n1695 = ( ~n21 & n1671 ) | ( ~n21 & n1694 ) | ( n1671 & n1694 ) ;
  assign n1696 = ( x0 & x3 ) | ( x0 & n689 ) | ( x3 & n689 ) ;
  assign n1697 = ( x0 & x3 ) | ( x0 & ~n689 ) | ( x3 & ~n689 ) ;
  assign n1698 = ( x4 & ~x8 ) | ( x4 & n1697 ) | ( ~x8 & n1697 ) ;
  assign n1699 = ~n1696 & n1698 ;
  assign n1700 = ~x3 & n145 ;
  assign n1701 = ( x0 & ~x4 ) | ( x0 & n1700 ) | ( ~x4 & n1700 ) ;
  assign n1702 = ~x0 & n1701 ;
  assign n1703 = x7 | n1702 ;
  assign n1704 = ( n1699 & n1702 ) | ( n1699 & n1703 ) | ( n1702 & n1703 ) ;
  assign n1705 = x1 | n1704 ;
  assign n1706 = x3 & x7 ;
  assign n1707 = x3 & ~n85 ;
  assign n1708 = ( n83 & n1706 ) | ( n83 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1709 = ~x0 & n1708 ;
  assign n1710 = x1 & ~n1709 ;
  assign n1711 = n1705 & ~n1710 ;
  assign n1712 = x2 | n1711 ;
  assign n1713 = ( x1 & ~x4 ) | ( x1 & n68 ) | ( ~x4 & n68 ) ;
  assign n1714 = ( x4 & ~x7 ) | ( x4 & n68 ) | ( ~x7 & n68 ) ;
  assign n1715 = ( x1 & x8 ) | ( x1 & ~n1714 ) | ( x8 & ~n1714 ) ;
  assign n1716 = ~n1713 & n1715 ;
  assign n1717 = ( ~x4 & n145 ) | ( ~x4 & n1716 ) | ( n145 & n1716 ) ;
  assign n1718 = n121 & ~n1717 ;
  assign n1719 = ( n121 & n1716 ) | ( n121 & ~n1718 ) | ( n1716 & ~n1718 ) ;
  assign n1720 = ~x0 & n1719 ;
  assign n1721 = x2 & ~n1720 ;
  assign n1722 = n1712 & ~n1721 ;
  assign n1723 = x5 | n1722 ;
  assign n1724 = ( n10 & n306 ) | ( n10 & ~n1656 ) | ( n306 & ~n1656 ) ;
  assign n1725 = x2 & ~n105 ;
  assign n1726 = n1724 & n1725 ;
  assign n1727 = ~x3 & n10 ;
  assign n1728 = ( ~n105 & n1725 ) | ( ~n105 & n1727 ) | ( n1725 & n1727 ) ;
  assign n1729 = ( x1 & n1726 ) | ( x1 & n1728 ) | ( n1726 & n1728 ) ;
  assign n1730 = n1725 & n1727 ;
  assign n1731 = x3 & n145 ;
  assign n1732 = ( ~n105 & n1725 ) | ( ~n105 & n1731 ) | ( n1725 & n1731 ) ;
  assign n1733 = ( x1 & n1730 ) | ( x1 & n1732 ) | ( n1730 & n1732 ) ;
  assign n1734 = x4 & ~n1733 ;
  assign n1735 = ( n1729 & n1733 ) | ( n1729 & ~n1734 ) | ( n1733 & ~n1734 ) ;
  assign n1736 = ~x0 & n1735 ;
  assign n1737 = x5 & ~n1736 ;
  assign n1738 = n1723 & ~n1737 ;
  assign n1739 = ~n20 & n463 ;
  assign n1740 = ( x4 & ~x7 ) | ( x4 & n721 ) | ( ~x7 & n721 ) ;
  assign n1741 = x4 & ~n1740 ;
  assign n1742 = n1740 | n1741 ;
  assign n1743 = ( ~x4 & n1741 ) | ( ~x4 & n1742 ) | ( n1741 & n1742 ) ;
  assign n1744 = ~x1 & n1743 ;
  assign n1745 = ~x1 & x7 ;
  assign n1746 = ( ~x2 & x4 ) | ( ~x2 & x8 ) | ( x4 & x8 ) ;
  assign n1747 = x2 & n1746 ;
  assign n1748 = ( ~n187 & n1746 ) | ( ~n187 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1749 = ( ~x1 & x7 ) | ( ~x1 & n1748 ) | ( x7 & n1748 ) ;
  assign n1750 = ( n1744 & ~n1745 ) | ( n1744 & n1749 ) | ( ~n1745 & n1749 ) ;
  assign n1751 = x3 & n1750 ;
  assign n1752 = ( x1 & ~x4 ) | ( x1 & x7 ) | ( ~x4 & x7 ) ;
  assign n1753 = ( x4 & ~x8 ) | ( x4 & n1752 ) | ( ~x8 & n1752 ) ;
  assign n1754 = ( x1 & x7 ) | ( x1 & n1753 ) | ( x7 & n1753 ) ;
  assign n1755 = n1752 & ~n1754 ;
  assign n1756 = ( n1753 & ~n1754 ) | ( n1753 & n1755 ) | ( ~n1754 & n1755 ) ;
  assign n1757 = x2 & ~n1756 ;
  assign n1758 = x1 & n145 ;
  assign n1759 = x2 | n1758 ;
  assign n1760 = ~n1757 & n1759 ;
  assign n1761 = x3 | n1760 ;
  assign n1762 = ( ~x3 & n1751 ) | ( ~x3 & n1761 ) | ( n1751 & n1761 ) ;
  assign n1763 = x6 & n1762 ;
  assign n1764 = x2 & n1563 ;
  assign n1765 = x3 | n1563 ;
  assign n1766 = ( x2 & ~x4 ) | ( x2 & n1765 ) | ( ~x4 & n1765 ) ;
  assign n1767 = ~n1764 & n1766 ;
  assign n1768 = ( x1 & ~x8 ) | ( x1 & n1767 ) | ( ~x8 & n1767 ) ;
  assign n1769 = ~x7 & n36 ;
  assign n1770 = ( x3 & x4 ) | ( x3 & ~n36 ) | ( x4 & ~n36 ) ;
  assign n1771 = ( x7 & n192 ) | ( x7 & ~n1770 ) | ( n192 & ~n1770 ) ;
  assign n1772 = ( x7 & n1769 ) | ( x7 & ~n1771 ) | ( n1769 & ~n1771 ) ;
  assign n1773 = ( x1 & x8 ) | ( x1 & ~n1772 ) | ( x8 & ~n1772 ) ;
  assign n1774 = n1768 & ~n1773 ;
  assign n1775 = ( x1 & ~n145 ) | ( x1 & n817 ) | ( ~n145 & n817 ) ;
  assign n1776 = n145 & n1775 ;
  assign n1777 = n1774 | n1776 ;
  assign n1778 = ~x6 & n1777 ;
  assign n1779 = n1763 | n1778 ;
  assign n1780 = ~x0 & n1779 ;
  assign n1781 = n99 | n1780 ;
  assign n1782 = ( n1739 & n1780 ) | ( n1739 & n1781 ) | ( n1780 & n1781 ) ;
  assign n1783 = x5 & ~n1782 ;
  assign n1784 = ( x2 & ~x7 ) | ( x2 & x8 ) | ( ~x7 & x8 ) ;
  assign n1785 = ( ~x2 & x4 ) | ( ~x2 & n1784 ) | ( x4 & n1784 ) ;
  assign n1786 = ( x4 & x8 ) | ( x4 & ~n1784 ) | ( x8 & ~n1784 ) ;
  assign n1787 = n1785 & ~n1786 ;
  assign n1788 = ( x1 & x6 ) | ( x1 & ~n1787 ) | ( x6 & ~n1787 ) ;
  assign n1789 = x4 & n57 ;
  assign n1790 = n68 & n1789 ;
  assign n1791 = x6 & n1790 ;
  assign n1792 = ( n1787 & n1788 ) | ( n1787 & n1791 ) | ( n1788 & n1791 ) ;
  assign n1793 = ( x1 & x4 ) | ( x1 & x6 ) | ( x4 & x6 ) ;
  assign n1794 = ( x2 & x7 ) | ( x2 & x8 ) | ( x7 & x8 ) ;
  assign n1795 = ( ~x3 & x8 ) | ( ~x3 & n1794 ) | ( x8 & n1794 ) ;
  assign n1796 = x8 & ~n1795 ;
  assign n1797 = n1795 | n1796 ;
  assign n1798 = ( ~x8 & n1796 ) | ( ~x8 & n1797 ) | ( n1796 & n1797 ) ;
  assign n1799 = x1 | x4 ;
  assign n1800 = ( x6 & n1798 ) | ( x6 & n1799 ) | ( n1798 & n1799 ) ;
  assign n1801 = ~n1793 & n1800 ;
  assign n1802 = ( ~x3 & n1792 ) | ( ~x3 & n1801 ) | ( n1792 & n1801 ) ;
  assign n1803 = ~x2 & x7 ;
  assign n1804 = ( x2 & x6 ) | ( x2 & n1803 ) | ( x6 & n1803 ) ;
  assign n1805 = ( x1 & x6 ) | ( x1 & n1803 ) | ( x6 & n1803 ) ;
  assign n1806 = ( n511 & n1804 ) | ( n511 & ~n1805 ) | ( n1804 & ~n1805 ) ;
  assign n1807 = x8 & ~n1806 ;
  assign n1808 = ~x1 & x6 ;
  assign n1809 = x1 & n597 ;
  assign n1810 = ( x1 & n1808 ) | ( x1 & ~n1809 ) | ( n1808 & ~n1809 ) ;
  assign n1811 = x2 & ~n1810 ;
  assign n1812 = x8 | n1811 ;
  assign n1813 = ~n1807 & n1812 ;
  assign n1814 = x4 & ~n1813 ;
  assign n1815 = ( x6 & ~x8 ) | ( x6 & n84 ) | ( ~x8 & n84 ) ;
  assign n1816 = ( ~x1 & x8 ) | ( ~x1 & n1815 ) | ( x8 & n1815 ) ;
  assign n1817 = ( x6 & x7 ) | ( x6 & ~n1816 ) | ( x7 & ~n1816 ) ;
  assign n1818 = ~n1815 & n1817 ;
  assign n1819 = x2 & n1818 ;
  assign n1820 = x4 | n1819 ;
  assign n1821 = ~n1814 & n1820 ;
  assign n1822 = ( x3 & n1801 ) | ( x3 & n1821 ) | ( n1801 & n1821 ) ;
  assign n1823 = n1802 | n1822 ;
  assign n1824 = ~x0 & n1823 ;
  assign n1825 = x5 | n1824 ;
  assign n1826 = ~n1783 & n1825 ;
  assign n1827 = n36 & n118 ;
  assign n1828 = ( x1 & n572 ) | ( x1 & n1827 ) | ( n572 & n1827 ) ;
  assign n1829 = ~x1 & n1828 ;
  assign n1830 = ( x2 & x6 ) | ( x2 & n83 ) | ( x6 & n83 ) ;
  assign n1831 = ~x2 & n1830 ;
  assign n1832 = ( x1 & ~x3 ) | ( x1 & n1831 ) | ( ~x3 & n1831 ) ;
  assign n1833 = ( x1 & x4 ) | ( x1 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n1834 = ( x1 & ~x7 ) | ( x1 & n1833 ) | ( ~x7 & n1833 ) ;
  assign n1835 = x1 & ~n1834 ;
  assign n1836 = n1834 | n1835 ;
  assign n1837 = ( ~x1 & n1835 ) | ( ~x1 & n1836 ) | ( n1835 & n1836 ) ;
  assign n1838 = ( ~x2 & x6 ) | ( ~x2 & n1837 ) | ( x6 & n1837 ) ;
  assign n1839 = ( ~x4 & x5 ) | ( ~x4 & x7 ) | ( x5 & x7 ) ;
  assign n1840 = ~x5 & n1839 ;
  assign n1841 = ( x4 & n1839 ) | ( x4 & n1840 ) | ( n1839 & n1840 ) ;
  assign n1842 = ~x1 & n1841 ;
  assign n1843 = ~x2 & n1842 ;
  assign n1844 = ~x6 & n1843 ;
  assign n1845 = ( n1837 & ~n1838 ) | ( n1837 & n1844 ) | ( ~n1838 & n1844 ) ;
  assign n1846 = ~x3 & n1845 ;
  assign n1847 = ( ~x1 & n1832 ) | ( ~x1 & n1846 ) | ( n1832 & n1846 ) ;
  assign n1848 = n99 & n551 ;
  assign n1849 = n22 & n1848 ;
  assign n1850 = ( ~n1829 & n1847 ) | ( ~n1829 & n1849 ) | ( n1847 & n1849 ) ;
  assign n1851 = x0 & ~n1849 ;
  assign n1852 = ( n1829 & n1850 ) | ( n1829 & ~n1851 ) | ( n1850 & ~n1851 ) ;
  assign n1853 = n1826 | n1852 ;
  assign n1854 = ( ~n1695 & n1738 ) | ( ~n1695 & n1853 ) | ( n1738 & n1853 ) ;
  assign n1855 = n1695 | n1854 ;
  assign n1856 = x1 & ~x5 ;
  assign n1857 = ( ~x0 & x3 ) | ( ~x0 & n1856 ) | ( x3 & n1856 ) ;
  assign n1858 = ( x1 & x3 ) | ( x1 & ~n1856 ) | ( x3 & ~n1856 ) ;
  assign n1859 = ( x5 & n1857 ) | ( x5 & ~n1858 ) | ( n1857 & ~n1858 ) ;
  assign n1860 = ( x1 & ~x7 ) | ( x1 & n120 ) | ( ~x7 & n120 ) ;
  assign n1861 = ~x1 & n1860 ;
  assign n1862 = x7 | n1861 ;
  assign n1863 = ( n1859 & n1861 ) | ( n1859 & n1862 ) | ( n1861 & n1862 ) ;
  assign n1864 = x2 | n1863 ;
  assign n1865 = ( ~x1 & x5 ) | ( ~x1 & n1706 ) | ( x5 & n1706 ) ;
  assign n1866 = ( x1 & ~x3 ) | ( x1 & n1706 ) | ( ~x3 & n1706 ) ;
  assign n1867 = ( x5 & x7 ) | ( x5 & ~n1866 ) | ( x7 & ~n1866 ) ;
  assign n1868 = ~n1865 & n1867 ;
  assign n1869 = ~x0 & n1868 ;
  assign n1870 = x2 & ~n1869 ;
  assign n1871 = n1864 & ~n1870 ;
  assign n1872 = ( n85 & ~n463 ) | ( n85 & n729 ) | ( ~n463 & n729 ) ;
  assign n1873 = n1871 & ~n1872 ;
  assign n1874 = ( x1 & x3 ) | ( x1 & ~x7 ) | ( x3 & ~x7 ) ;
  assign n1875 = n949 & ~n1874 ;
  assign n1876 = x0 | n1875 ;
  assign n1877 = x4 | n1575 ;
  assign n1878 = x1 | n1877 ;
  assign n1879 = x0 & n1878 ;
  assign n1880 = n1876 & ~n1879 ;
  assign n1881 = n1156 & n1880 ;
  assign n1882 = n52 & n98 ;
  assign n1883 = ( n26 & ~n145 ) | ( n26 & n1882 ) | ( ~n145 & n1882 ) ;
  assign n1884 = n145 & n1883 ;
  assign n1885 = ( ~x3 & x7 ) | ( ~x3 & x8 ) | ( x7 & x8 ) ;
  assign n1886 = ( x3 & ~x8 ) | ( x3 & n1885 ) | ( ~x8 & n1885 ) ;
  assign n1887 = ~x6 & n1885 ;
  assign n1888 = ( ~x7 & n1885 ) | ( ~x7 & n1887 ) | ( n1885 & n1887 ) ;
  assign n1889 = n1886 | n1888 ;
  assign n1890 = x1 & n1889 ;
  assign n1891 = x3 | n58 ;
  assign n1892 = ~x1 & n1891 ;
  assign n1893 = n1890 | n1892 ;
  assign n1894 = x4 & ~n1893 ;
  assign n1895 = ~x1 & x8 ;
  assign n1896 = ( x6 & n306 ) | ( x6 & n1895 ) | ( n306 & n1895 ) ;
  assign n1897 = ( x3 & ~x6 ) | ( x3 & n1896 ) | ( ~x6 & n1896 ) ;
  assign n1898 = ( ~x8 & n1895 ) | ( ~x8 & n1897 ) | ( n1895 & n1897 ) ;
  assign n1899 = ( ~n1895 & n1896 ) | ( ~n1895 & n1898 ) | ( n1896 & n1898 ) ;
  assign n1900 = ~n58 & n121 ;
  assign n1901 = x7 | n1900 ;
  assign n1902 = ( n1899 & n1900 ) | ( n1899 & n1901 ) | ( n1900 & n1901 ) ;
  assign n1903 = x4 | n1902 ;
  assign n1904 = ( ~x4 & n1894 ) | ( ~x4 & n1903 ) | ( n1894 & n1903 ) ;
  assign n1905 = ( ~x0 & x5 ) | ( ~x0 & n1904 ) | ( x5 & n1904 ) ;
  assign n1906 = x7 & ~n880 ;
  assign n1907 = ~x6 & n1906 ;
  assign n1908 = ~x3 & n1907 ;
  assign n1909 = x6 & n26 ;
  assign n1910 = ~n20 & n1909 ;
  assign n1911 = ( x3 & ~x4 ) | ( x3 & x8 ) | ( ~x4 & x8 ) ;
  assign n1912 = ( ~x3 & x7 ) | ( ~x3 & n1911 ) | ( x7 & n1911 ) ;
  assign n1913 = ( ~x4 & x8 ) | ( ~x4 & n1912 ) | ( x8 & n1912 ) ;
  assign n1914 = ~n1911 & n1913 ;
  assign n1915 = ( ~n1912 & n1913 ) | ( ~n1912 & n1914 ) | ( n1913 & n1914 ) ;
  assign n1916 = n1910 | n1915 ;
  assign n1917 = ( n1907 & ~n1908 ) | ( n1907 & n1916 ) | ( ~n1908 & n1916 ) ;
  assign n1918 = x1 | n1917 ;
  assign n1919 = x3 & ~x8 ;
  assign n1920 = ( x3 & ~x7 ) | ( x3 & n347 ) | ( ~x7 & n347 ) ;
  assign n1921 = n347 | n1920 ;
  assign n1922 = ~n1919 & n1921 ;
  assign n1923 = ~x6 & n1922 ;
  assign n1924 = x1 & ~n1923 ;
  assign n1925 = n1918 & ~n1924 ;
  assign n1926 = ( x6 & ~x8 ) | ( x6 & n1146 ) | ( ~x8 & n1146 ) ;
  assign n1927 = x8 & n1926 ;
  assign n1928 = n1926 & ~n1927 ;
  assign n1929 = ( x8 & ~n1927 ) | ( x8 & n1928 ) | ( ~n1927 & n1928 ) ;
  assign n1930 = ( x3 & ~x4 ) | ( x3 & n1929 ) | ( ~x4 & n1929 ) ;
  assign n1931 = ( n26 & ~n1925 ) | ( n26 & n1930 ) | ( ~n1925 & n1930 ) ;
  assign n1932 = ( x0 & x5 ) | ( x0 & n1931 ) | ( x5 & n1931 ) ;
  assign n1933 = n1905 & ~n1932 ;
  assign n1934 = n1884 | n1933 ;
  assign n1935 = ( n1880 & ~n1881 ) | ( n1880 & n1934 ) | ( ~n1881 & n1934 ) ;
  assign n1936 = x2 | n1935 ;
  assign n1937 = ( ~x3 & x8 ) | ( ~x3 & n232 ) | ( x8 & n232 ) ;
  assign n1938 = ( x5 & x7 ) | ( x5 & n1937 ) | ( x7 & n1937 ) ;
  assign n1939 = ~n232 & n1938 ;
  assign n1940 = ( ~n1937 & n1938 ) | ( ~n1937 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1941 = x1 | n1940 ;
  assign n1942 = x3 | n134 ;
  assign n1943 = x1 & n1942 ;
  assign n1944 = n1941 & ~n1943 ;
  assign n1945 = x4 & n1944 ;
  assign n1946 = ( ~x3 & x5 ) | ( ~x3 & x7 ) | ( x5 & x7 ) ;
  assign n1947 = ( x1 & x5 ) | ( x1 & ~n1946 ) | ( x5 & ~n1946 ) ;
  assign n1948 = ( ~x5 & x7 ) | ( ~x5 & n1947 ) | ( x7 & n1947 ) ;
  assign n1949 = n1946 & n1948 ;
  assign n1950 = x1 & ~n1949 ;
  assign n1951 = ( n1947 & n1949 ) | ( n1947 & ~n1950 ) | ( n1949 & ~n1950 ) ;
  assign n1952 = x8 & n1951 ;
  assign n1953 = ( x1 & ~x3 ) | ( x1 & x7 ) | ( ~x3 & x7 ) ;
  assign n1954 = ( ~x1 & x3 ) | ( ~x1 & x8 ) | ( x3 & x8 ) ;
  assign n1955 = n1953 | n1954 ;
  assign n1956 = ~n1952 & n1955 ;
  assign n1957 = ( x5 & n1952 ) | ( x5 & ~n1956 ) | ( n1952 & ~n1956 ) ;
  assign n1958 = x4 | n1957 ;
  assign n1959 = ( ~x4 & n1945 ) | ( ~x4 & n1958 ) | ( n1945 & n1958 ) ;
  assign n1960 = x6 & ~n1959 ;
  assign n1961 = x1 & x5 ;
  assign n1962 = x3 & x5 ;
  assign n1963 = ( x1 & ~x7 ) | ( x1 & n1962 ) | ( ~x7 & n1962 ) ;
  assign n1964 = ( n738 & ~n1961 ) | ( n738 & n1963 ) | ( ~n1961 & n1963 ) ;
  assign n1965 = x4 & n1964 ;
  assign n1966 = ( x4 & ~x7 ) | ( x4 & n1513 ) | ( ~x7 & n1513 ) ;
  assign n1967 = ( ~n83 & n1965 ) | ( ~n83 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1968 = x8 & n1967 ;
  assign n1969 = x6 | n1968 ;
  assign n1970 = ~n1960 & n1969 ;
  assign n1971 = ( ~x1 & x8 ) | ( ~x1 & n394 ) | ( x8 & n394 ) ;
  assign n1972 = ( x7 & x8 ) | ( x7 & ~n394 ) | ( x8 & ~n394 ) ;
  assign n1973 = ( ~x1 & x4 ) | ( ~x1 & n1972 ) | ( x4 & n1972 ) ;
  assign n1974 = ~n1971 & n1973 ;
  assign n1975 = x5 & ~n1974 ;
  assign n1976 = n10 & ~n1799 ;
  assign n1977 = x5 | n1976 ;
  assign n1978 = ~n1975 & n1977 ;
  assign n1979 = ( ~x3 & x6 ) | ( ~x3 & n1978 ) | ( x6 & n1978 ) ;
  assign n1980 = ( ~n1465 & n1970 ) | ( ~n1465 & n1979 ) | ( n1970 & n1979 ) ;
  assign n1981 = ~x0 & n1980 ;
  assign n1982 = x2 & ~n1981 ;
  assign n1983 = n1936 & ~n1982 ;
  assign n1984 = ( ~x3 & x4 ) | ( ~x3 & x7 ) | ( x4 & x7 ) ;
  assign n1985 = ( x1 & x3 ) | ( x1 & n1984 ) | ( x3 & n1984 ) ;
  assign n1986 = ( x3 & x7 ) | ( x3 & ~n1985 ) | ( x7 & ~n1985 ) ;
  assign n1987 = n1984 & n1986 ;
  assign n1988 = ( x1 & ~n1985 ) | ( x1 & n1987 ) | ( ~n1985 & n1987 ) ;
  assign n1989 = x2 & ~n1988 ;
  assign n1990 = x3 & ~n346 ;
  assign n1991 = ( x4 & ~n346 ) | ( x4 & n1990 ) | ( ~n346 & n1990 ) ;
  assign n1992 = x1 & n1991 ;
  assign n1993 = x2 | n1992 ;
  assign n1994 = ~n1989 & n1993 ;
  assign n1995 = x6 & ~n1994 ;
  assign n1996 = ( x1 & x3 ) | ( x1 & ~n1328 ) | ( x3 & ~n1328 ) ;
  assign n1997 = ( x2 & x4 ) | ( x2 & ~n1996 ) | ( x4 & ~n1996 ) ;
  assign n1998 = ~n1328 & n1997 ;
  assign n1999 = ( n1996 & n1997 ) | ( n1996 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2000 = ~x7 & n1999 ;
  assign n2001 = x6 | n2000 ;
  assign n2002 = ~n1995 & n2001 ;
  assign n2003 = x0 | n2002 ;
  assign n2004 = n26 & ~n566 ;
  assign n2005 = ~n15 & n2004 ;
  assign n2006 = x0 & ~n2005 ;
  assign n2007 = n2003 & ~n2006 ;
  assign n2008 = x5 & n2007 ;
  assign n2009 = ( x2 & ~x3 ) | ( x2 & x6 ) | ( ~x3 & x6 ) ;
  assign n2010 = x6 & ~n2009 ;
  assign n2011 = ( x1 & x2 ) | ( x1 & n2010 ) | ( x2 & n2010 ) ;
  assign n2012 = ( ~n2009 & n2010 ) | ( ~n2009 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = ( x0 & ~n243 ) | ( x0 & n2012 ) | ( ~n243 & n2012 ) ;
  assign n2014 = ( x2 & n98 ) | ( x2 & n1465 ) | ( n98 & n1465 ) ;
  assign n2015 = ~x2 & n2014 ;
  assign n2016 = ~n243 & n2015 ;
  assign n2017 = ( ~x0 & n2013 ) | ( ~x0 & n2016 ) | ( n2013 & n2016 ) ;
  assign n2018 = ~x6 & n26 ;
  assign n2019 = n320 & ~n2018 ;
  assign n2020 = ( x4 & n106 ) | ( x4 & n1420 ) | ( n106 & n1420 ) ;
  assign n2021 = ~x4 & n2020 ;
  assign n2022 = ( x1 & x7 ) | ( x1 & ~n1420 ) | ( x7 & ~n1420 ) ;
  assign n2023 = ( ~x1 & x3 ) | ( ~x1 & n2022 ) | ( x3 & n2022 ) ;
  assign n2024 = ( x6 & ~x7 ) | ( x6 & n2023 ) | ( ~x7 & n2023 ) ;
  assign n2025 = n2022 & n2024 ;
  assign n2026 = ~x1 & n1114 ;
  assign n2027 = x4 & ~n2026 ;
  assign n2028 = ( n2025 & n2026 ) | ( n2025 & ~n2027 ) | ( n2026 & ~n2027 ) ;
  assign n2029 = ( ~x0 & x2 ) | ( ~x0 & n2028 ) | ( x2 & n2028 ) ;
  assign n2030 = ( x1 & x7 ) | ( x1 & ~n1575 ) | ( x7 & ~n1575 ) ;
  assign n2031 = ( x1 & x6 ) | ( x1 & ~n1575 ) | ( x6 & ~n1575 ) ;
  assign n2032 = ( n597 & n2030 ) | ( n597 & ~n2031 ) | ( n2030 & ~n2031 ) ;
  assign n2033 = x4 | n2032 ;
  assign n2034 = n121 & n551 ;
  assign n2035 = x4 & ~n2034 ;
  assign n2036 = n2033 & ~n2035 ;
  assign n2037 = ( x0 & x2 ) | ( x0 & ~n2036 ) | ( x2 & ~n2036 ) ;
  assign n2038 = n2029 & ~n2037 ;
  assign n2039 = n2021 | n2038 ;
  assign n2040 = ( n320 & ~n2019 ) | ( n320 & n2039 ) | ( ~n2019 & n2039 ) ;
  assign n2041 = n2017 | n2040 ;
  assign n2042 = ~x5 & n2041 ;
  assign n2043 = n2008 | n2042 ;
  assign n2044 = n1983 | n2043 ;
  assign n2045 = ( n1871 & ~n1873 ) | ( n1871 & n2044 ) | ( ~n1873 & n2044 ) ;
  assign n2046 = ( x3 & ~x5 ) | ( x3 & x6 ) | ( ~x5 & x6 ) ;
  assign n2047 = ( x4 & ~x6 ) | ( x4 & n2046 ) | ( ~x6 & n2046 ) ;
  assign n2048 = ( x3 & x4 ) | ( x3 & ~n2046 ) | ( x4 & ~n2046 ) ;
  assign n2049 = n2047 & ~n2048 ;
  assign n2050 = ( x0 & ~x1 ) | ( x0 & n2049 ) | ( ~x1 & n2049 ) ;
  assign n2051 = n1278 & ~n1356 ;
  assign n2052 = ~x0 & n2051 ;
  assign n2053 = ( n2049 & ~n2050 ) | ( n2049 & n2052 ) | ( ~n2050 & n2052 ) ;
  assign n2054 = ( x3 & x5 ) | ( x3 & x6 ) | ( x5 & x6 ) ;
  assign n2055 = ( ~x4 & x6 ) | ( ~x4 & n2054 ) | ( x6 & n2054 ) ;
  assign n2056 = x6 & ~n2055 ;
  assign n2057 = n2055 | n2056 ;
  assign n2058 = ( ~x6 & n2056 ) | ( ~x6 & n2057 ) | ( n2056 & n2057 ) ;
  assign n2059 = ( x1 & n1259 ) | ( x1 & ~n2058 ) | ( n1259 & ~n2058 ) ;
  assign n2060 = n2058 & n2059 ;
  assign n2061 = ( n1359 & ~n2053 ) | ( n1359 & n2060 ) | ( ~n2053 & n2060 ) ;
  assign n2062 = x2 & ~n2060 ;
  assign n2063 = ( n2053 & n2061 ) | ( n2053 & ~n2062 ) | ( n2061 & ~n2062 ) ;
  assign n2064 = ~n21 & n2063 ;
  assign n2065 = ( x5 & x8 ) | ( x5 & ~n378 ) | ( x8 & ~n378 ) ;
  assign n2066 = ( ~x0 & x5 ) | ( ~x0 & n378 ) | ( x5 & n378 ) ;
  assign n2067 = ( ~x2 & x8 ) | ( ~x2 & n2066 ) | ( x8 & n2066 ) ;
  assign n2068 = n2065 & ~n2067 ;
  assign n2069 = ~x7 & n2068 ;
  assign n2070 = ( ~x5 & n589 ) | ( ~x5 & n1803 ) | ( n589 & n1803 ) ;
  assign n2071 = n2069 | n2070 ;
  assign n2072 = ( x0 & n2069 ) | ( x0 & n2071 ) | ( n2069 & n2071 ) ;
  assign n2073 = x4 & ~n2072 ;
  assign n2074 = ~x7 & n1238 ;
  assign n2075 = ( x2 & x5 ) | ( x2 & ~n2074 ) | ( x5 & ~n2074 ) ;
  assign n2076 = ( n1238 & n2074 ) | ( n1238 & ~n2075 ) | ( n2074 & ~n2075 ) ;
  assign n2077 = ~x0 & n2076 ;
  assign n2078 = x4 | n2077 ;
  assign n2079 = ~n2073 & n2078 ;
  assign n2080 = x1 & n2079 ;
  assign n2081 = ( n145 & n171 ) | ( n145 & n770 ) | ( n171 & n770 ) ;
  assign n2082 = ( ~x8 & n145 ) | ( ~x8 & n2081 ) | ( n145 & n2081 ) ;
  assign n2083 = ( x4 & ~n101 ) | ( x4 & n2082 ) | ( ~n101 & n2082 ) ;
  assign n2084 = n2082 & ~n2083 ;
  assign n2085 = ( x1 & n812 ) | ( x1 & n880 ) | ( n812 & n880 ) ;
  assign n2086 = ~n880 & n2085 ;
  assign n2087 = ( ~x4 & n695 ) | ( ~x4 & n2086 ) | ( n695 & n2086 ) ;
  assign n2088 = n57 & ~n2087 ;
  assign n2089 = ( n57 & n2086 ) | ( n57 & ~n2088 ) | ( n2086 & ~n2088 ) ;
  assign n2090 = x0 | n2089 ;
  assign n2091 = n15 | n1537 ;
  assign n2092 = x0 & n2091 ;
  assign n2093 = n2090 & ~n2092 ;
  assign n2094 = n2084 | n2093 ;
  assign n2095 = ( n2079 & ~n2080 ) | ( n2079 & n2094 ) | ( ~n2080 & n2094 ) ;
  assign n2096 = x3 | n2095 ;
  assign n2097 = ( x5 & ~x7 ) | ( x5 & n155 ) | ( ~x7 & n155 ) ;
  assign n2098 = ( x7 & x8 ) | ( x7 & ~n155 ) | ( x8 & ~n155 ) ;
  assign n2099 = ( ~n38 & n2097 ) | ( ~n38 & n2098 ) | ( n2097 & n2098 ) ;
  assign n2100 = x4 & ~n2099 ;
  assign n2101 = x2 & n68 ;
  assign n2102 = x4 | n2101 ;
  assign n2103 = ~n2100 & n2102 ;
  assign n2104 = x1 & n2103 ;
  assign n2105 = ( x5 & n312 ) | ( x5 & ~n1803 ) | ( n312 & ~n1803 ) ;
  assign n2106 = ( ~x5 & x7 ) | ( ~x5 & n2105 ) | ( x7 & n2105 ) ;
  assign n2107 = ( ~x2 & n312 ) | ( ~x2 & n2106 ) | ( n312 & n2106 ) ;
  assign n2108 = ( ~n312 & n2105 ) | ( ~n312 & n2107 ) | ( n2105 & n2107 ) ;
  assign n2109 = ~x4 & n2108 ;
  assign n2110 = ~x2 & n247 ;
  assign n2111 = x4 & ~n2110 ;
  assign n2112 = n2109 | n2111 ;
  assign n2113 = ~x1 & n2112 ;
  assign n2114 = ( x1 & ~n2104 ) | ( x1 & n2113 ) | ( ~n2104 & n2113 ) ;
  assign n2115 = x0 | n2114 ;
  assign n2116 = x3 & n2115 ;
  assign n2117 = n2096 & ~n2116 ;
  assign n2118 = ( x2 & ~x3 ) | ( x2 & n921 ) | ( ~x3 & n921 ) ;
  assign n2119 = x2 | n2118 ;
  assign n2120 = x2 & n2118 ;
  assign n2121 = n2119 & ~n2120 ;
  assign n2122 = ( x0 & ~x7 ) | ( x0 & n2121 ) | ( ~x7 & n2121 ) ;
  assign n2123 = ~n15 & n1114 ;
  assign n2124 = ~x0 & n2123 ;
  assign n2125 = ( n2121 & ~n2122 ) | ( n2121 & n2124 ) | ( ~n2122 & n2124 ) ;
  assign n2126 = ( x3 & n320 ) | ( x3 & n785 ) | ( n320 & n785 ) ;
  assign n2127 = ~x3 & n2126 ;
  assign n2128 = n144 & ~n811 ;
  assign n2129 = ( x5 & x7 ) | ( x5 & n1106 ) | ( x7 & n1106 ) ;
  assign n2130 = ( x4 & x7 ) | ( x4 & ~n2129 ) | ( x7 & ~n2129 ) ;
  assign n2131 = n1106 | n2130 ;
  assign n2132 = ( x5 & ~n2129 ) | ( x5 & n2131 ) | ( ~n2129 & n2131 ) ;
  assign n2133 = x6 & ~n2132 ;
  assign n2134 = ~x2 & n2133 ;
  assign n2135 = ( x2 & ~x7 ) | ( x2 & n1398 ) | ( ~x7 & n1398 ) ;
  assign n2136 = x2 & ~n2135 ;
  assign n2137 = n2135 | n2136 ;
  assign n2138 = ( ~x2 & n2136 ) | ( ~x2 & n2137 ) | ( n2136 & n2137 ) ;
  assign n2139 = ~x2 & n2018 ;
  assign n2140 = x6 | n2139 ;
  assign n2141 = ( n2138 & n2139 ) | ( n2138 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = n2134 | n2141 ;
  assign n2143 = ( n144 & ~n2128 ) | ( n144 & n2142 ) | ( ~n2128 & n2142 ) ;
  assign n2144 = ( ~x0 & x1 ) | ( ~x0 & n2143 ) | ( x1 & n2143 ) ;
  assign n2145 = ( ~x3 & x6 ) | ( ~x3 & x7 ) | ( x6 & x7 ) ;
  assign n2146 = x7 & n2145 ;
  assign n2147 = ( ~x3 & x4 ) | ( ~x3 & n2146 ) | ( x4 & n2146 ) ;
  assign n2148 = ( n330 & n2145 ) | ( n330 & ~n2147 ) | ( n2145 & ~n2147 ) ;
  assign n2149 = x5 | n2148 ;
  assign n2150 = n60 & ~n566 ;
  assign n2151 = x5 & ~n2150 ;
  assign n2152 = n2149 & ~n2151 ;
  assign n2153 = x2 | n2152 ;
  assign n2154 = n26 & n552 ;
  assign n2155 = x2 & ~n2154 ;
  assign n2156 = n2153 & ~n2155 ;
  assign n2157 = ( x0 & x1 ) | ( x0 & ~n2156 ) | ( x1 & ~n2156 ) ;
  assign n2158 = n2144 & ~n2157 ;
  assign n2159 = ( ~n2125 & n2127 ) | ( ~n2125 & n2158 ) | ( n2127 & n2158 ) ;
  assign n2160 = n1426 & ~n2158 ;
  assign n2161 = ( n2125 & n2159 ) | ( n2125 & ~n2160 ) | ( n2159 & ~n2160 ) ;
  assign n2162 = x8 & ~n2161 ;
  assign n2163 = x3 | n798 ;
  assign n2164 = x3 & n799 ;
  assign n2165 = n2163 & ~n2164 ;
  assign n2166 = x4 & ~n2165 ;
  assign n2167 = x3 & n171 ;
  assign n2168 = x4 | n2167 ;
  assign n2169 = ~n2166 & n2168 ;
  assign n2170 = ~x5 & n144 ;
  assign n2171 = n572 & n2170 ;
  assign n2172 = x6 & ~n2171 ;
  assign n2173 = ( n2169 & n2171 ) | ( n2169 & ~n2172 ) | ( n2171 & ~n2172 ) ;
  assign n2174 = ( x3 & x4 ) | ( x3 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n2175 = ( x3 & ~x7 ) | ( x3 & n2174 ) | ( ~x7 & n2174 ) ;
  assign n2176 = x3 & ~n2175 ;
  assign n2177 = n2175 | n2176 ;
  assign n2178 = ( ~x3 & n2176 ) | ( ~x3 & n2177 ) | ( n2176 & n2177 ) ;
  assign n2179 = ( x2 & x6 ) | ( x2 & n2178 ) | ( x6 & n2178 ) ;
  assign n2180 = ( x1 & ~x6 ) | ( x1 & n2179 ) | ( ~x6 & n2179 ) ;
  assign n2181 = ( x1 & x2 ) | ( x1 & ~n2179 ) | ( x2 & ~n2179 ) ;
  assign n2182 = n2180 & ~n2181 ;
  assign n2183 = ( ~x1 & n2173 ) | ( ~x1 & n2182 ) | ( n2173 & n2182 ) ;
  assign n2184 = x3 & ~x6 ;
  assign n2185 = ( ~x4 & x7 ) | ( ~x4 & n2184 ) | ( x7 & n2184 ) ;
  assign n2186 = ( x6 & ~x7 ) | ( x6 & n2184 ) | ( ~x7 & n2184 ) ;
  assign n2187 = ( ~x3 & x4 ) | ( ~x3 & n2186 ) | ( x4 & n2186 ) ;
  assign n2188 = n2185 | n2187 ;
  assign n2189 = x2 | n2188 ;
  assign n2190 = n430 & n551 ;
  assign n2191 = ( x2 & x3 ) | ( x2 & ~x6 ) | ( x3 & ~x6 ) ;
  assign n2192 = ( x2 & ~x7 ) | ( x2 & n2191 ) | ( ~x7 & n2191 ) ;
  assign n2193 = x2 & ~n2192 ;
  assign n2194 = n2192 | n2193 ;
  assign n2195 = ( ~x2 & n2193 ) | ( ~x2 & n2194 ) | ( n2193 & n2194 ) ;
  assign n2196 = n2190 | n2195 ;
  assign n2197 = ( ~n2188 & n2189 ) | ( ~n2188 & n2196 ) | ( n2189 & n2196 ) ;
  assign n2198 = x5 & ~n2197 ;
  assign n2199 = ( x7 & n53 ) | ( x7 & ~n1984 ) | ( n53 & ~n1984 ) ;
  assign n2200 = ( ~x2 & n1984 ) | ( ~x2 & n2199 ) | ( n1984 & n2199 ) ;
  assign n2201 = ( ~x7 & n2199 ) | ( ~x7 & n2200 ) | ( n2199 & n2200 ) ;
  assign n2202 = x6 | n2201 ;
  assign n2203 = ~x5 & n2202 ;
  assign n2204 = n2198 | n2203 ;
  assign n2205 = ( x1 & n2182 ) | ( x1 & ~n2204 ) | ( n2182 & ~n2204 ) ;
  assign n2206 = n2183 | n2205 ;
  assign n2207 = ~x0 & n2206 ;
  assign n2208 = x8 | n2207 ;
  assign n2209 = ~n2162 & n2208 ;
  assign n2210 = n2117 | n2209 ;
  assign n2211 = ( n2063 & ~n2064 ) | ( n2063 & n2210 ) | ( ~n2064 & n2210 ) ;
  assign n2212 = x0 & x3 ;
  assign n2213 = ( ~x4 & x5 ) | ( ~x4 & n2212 ) | ( x5 & n2212 ) ;
  assign n2214 = ( x3 & x5 ) | ( x3 & ~n2212 ) | ( x5 & ~n2212 ) ;
  assign n2215 = ( x0 & ~x4 ) | ( x0 & n2214 ) | ( ~x4 & n2214 ) ;
  assign n2216 = ~n2213 & n2215 ;
  assign n2217 = ( x1 & x2 ) | ( x1 & n2216 ) | ( x2 & n2216 ) ;
  assign n2218 = ( x4 & n101 ) | ( x4 & n672 ) | ( n101 & n672 ) ;
  assign n2219 = ~x4 & n2218 ;
  assign n2220 = ~x2 & n2219 ;
  assign n2221 = ( n2216 & ~n2217 ) | ( n2216 & n2220 ) | ( ~n2217 & n2220 ) ;
  assign n2222 = ( ~x3 & n67 ) | ( ~x3 & n2221 ) | ( n67 & n2221 ) ;
  assign n2223 = n106 & ~n2222 ;
  assign n2224 = ( n106 & n2221 ) | ( n106 & ~n2223 ) | ( n2221 & ~n2223 ) ;
  assign n2225 = n762 & n2224 ;
  assign n2226 = ( ~n576 & n613 ) | ( ~n576 & n1895 ) | ( n613 & n1895 ) ;
  assign n2227 = ( x3 & ~x7 ) | ( x3 & n2226 ) | ( ~x7 & n2226 ) ;
  assign n2228 = ~x3 & n2227 ;
  assign n2229 = ( x7 & n2227 ) | ( x7 & n2228 ) | ( n2227 & n2228 ) ;
  assign n2230 = n1356 & ~n2229 ;
  assign n2231 = ( n284 & n2229 ) | ( n284 & ~n2230 ) | ( n2229 & ~n2230 ) ;
  assign n2232 = x6 & ~n2231 ;
  assign n2233 = x5 & ~n1955 ;
  assign n2234 = x6 | n2233 ;
  assign n2235 = ~n2232 & n2234 ;
  assign n2236 = ~x2 & n2235 ;
  assign n2237 = ( x5 & ~x6 ) | ( x5 & x8 ) | ( ~x6 & x8 ) ;
  assign n2238 = ( x7 & x8 ) | ( x7 & ~n2237 ) | ( x8 & ~n2237 ) ;
  assign n2239 = ( ~x5 & x7 ) | ( ~x5 & n2237 ) | ( x7 & n2237 ) ;
  assign n2240 = n2238 & ~n2239 ;
  assign n2241 = ( ~x1 & x3 ) | ( ~x1 & n2240 ) | ( x3 & n2240 ) ;
  assign n2242 = x5 & n21 ;
  assign n2243 = ~x6 & n2242 ;
  assign n2244 = ( x1 & x3 ) | ( x1 & n2243 ) | ( x3 & n2243 ) ;
  assign n2245 = n2241 & n2244 ;
  assign n2246 = ~x1 & n884 ;
  assign n2247 = n37 & n2246 ;
  assign n2248 = n2245 | n2247 ;
  assign n2249 = x2 & n2248 ;
  assign n2250 = n2236 | n2249 ;
  assign n2251 = ( x2 & ~x6 ) | ( x2 & n832 ) | ( ~x6 & n832 ) ;
  assign n2252 = x2 & ~n2251 ;
  assign n2253 = n2251 | n2252 ;
  assign n2254 = ( ~x2 & n2252 ) | ( ~x2 & n2253 ) | ( n2252 & n2253 ) ;
  assign n2255 = ( x1 & n21 ) | ( x1 & n2254 ) | ( n21 & n2254 ) ;
  assign n2256 = ~x3 & n105 ;
  assign n2257 = n596 & n2256 ;
  assign n2258 = ~n21 & n2257 ;
  assign n2259 = ( n2254 & ~n2255 ) | ( n2254 & n2258 ) | ( ~n2255 & n2258 ) ;
  assign n2260 = ~x5 & n57 ;
  assign n2261 = x6 & ~n20 ;
  assign n2262 = n2260 & n2261 ;
  assign n2263 = ( x1 & ~x2 ) | ( x1 & n2262 ) | ( ~x2 & n2262 ) ;
  assign n2264 = n884 & ~n2263 ;
  assign n2265 = ( n884 & n2262 ) | ( n884 & ~n2264 ) | ( n2262 & ~n2264 ) ;
  assign n2266 = ( ~x0 & n2259 ) | ( ~x0 & n2265 ) | ( n2259 & n2265 ) ;
  assign n2267 = ~n2250 & n2266 ;
  assign n2268 = ( ~x0 & n2250 ) | ( ~x0 & n2267 ) | ( n2250 & n2267 ) ;
  assign n2269 = ( n99 & n145 ) | ( n99 & n2268 ) | ( n145 & n2268 ) ;
  assign n2270 = n52 & ~n2269 ;
  assign n2271 = ( n52 & n2268 ) | ( n52 & ~n2270 ) | ( n2268 & ~n2270 ) ;
  assign n2272 = ( x5 & ~x7 ) | ( x5 & n158 ) | ( ~x7 & n158 ) ;
  assign n2273 = x7 & n2272 ;
  assign n2274 = n2272 & ~n2273 ;
  assign n2275 = ( x7 & ~n2273 ) | ( x7 & n2274 ) | ( ~n2273 & n2274 ) ;
  assign n2276 = x4 & ~n2275 ;
  assign n2277 = x2 & n2276 ;
  assign n2278 = n811 | n2277 ;
  assign n2279 = ( ~n630 & n2277 ) | ( ~n630 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2280 = ( ~x0 & x1 ) | ( ~x0 & n2279 ) | ( x1 & n2279 ) ;
  assign n2281 = ( x5 & x7 ) | ( x5 & ~n1310 ) | ( x7 & ~n1310 ) ;
  assign n2282 = ( x4 & ~x6 ) | ( x4 & n2281 ) | ( ~x6 & n2281 ) ;
  assign n2283 = n1310 | n2282 ;
  assign n2284 = ( ~n2281 & n2282 ) | ( ~n2281 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2285 = x3 | n2284 ;
  assign n2286 = x2 | n2285 ;
  assign n2287 = ( x0 & x1 ) | ( x0 & n2286 ) | ( x1 & n2286 ) ;
  assign n2288 = n2280 & ~n2287 ;
  assign n2289 = ( n22 & n99 ) | ( n22 & n2288 ) | ( n99 & n2288 ) ;
  assign n2290 = n566 | n2289 ;
  assign n2291 = ( ~n566 & n2288 ) | ( ~n566 & n2290 ) | ( n2288 & n2290 ) ;
  assign n2292 = ( x4 & n2271 ) | ( x4 & n2291 ) | ( n2271 & n2291 ) ;
  assign n2293 = ( x6 & ~x8 ) | ( x6 & n1885 ) | ( ~x8 & n1885 ) ;
  assign n2294 = ( ~x7 & x8 ) | ( ~x7 & n2293 ) | ( x8 & n2293 ) ;
  assign n2295 = ~n1885 & n2294 ;
  assign n2296 = ( ~x6 & n2293 ) | ( ~x6 & n2295 ) | ( n2293 & n2295 ) ;
  assign n2297 = x1 | n2296 ;
  assign n2298 = ~x3 & n258 ;
  assign n2299 = x1 & ~n2298 ;
  assign n2300 = n2297 & ~n2299 ;
  assign n2301 = ( x7 & x8 ) | ( x7 & n122 ) | ( x8 & n122 ) ;
  assign n2302 = ( x6 & ~x7 ) | ( x6 & n2301 ) | ( ~x7 & n2301 ) ;
  assign n2303 = ( x6 & x8 ) | ( x6 & ~n2301 ) | ( x8 & ~n2301 ) ;
  assign n2304 = n2302 & ~n2303 ;
  assign n2305 = x0 & ~n2304 ;
  assign n2306 = ( n2300 & n2304 ) | ( n2300 & ~n2305 ) | ( n2304 & ~n2305 ) ;
  assign n2307 = x2 | n2306 ;
  assign n2308 = ~n74 & n584 ;
  assign n2309 = x3 | x8 ;
  assign n2310 = ( ~x1 & x3 ) | ( ~x1 & n1465 ) | ( x3 & n1465 ) ;
  assign n2311 = ( x1 & x8 ) | ( x1 & ~n1465 ) | ( x8 & ~n1465 ) ;
  assign n2312 = ( ~n2309 & n2310 ) | ( ~n2309 & n2311 ) | ( n2310 & n2311 ) ;
  assign n2313 = ~x7 & n2312 ;
  assign n2314 = ( ~x6 & n566 ) | ( ~x6 & n597 ) | ( n566 & n597 ) ;
  assign n2315 = ( x3 & x8 ) | ( x3 & ~n2314 ) | ( x8 & ~n2314 ) ;
  assign n2316 = ( x1 & ~x3 ) | ( x1 & n2315 ) | ( ~x3 & n2315 ) ;
  assign n2317 = ( x1 & x8 ) | ( x1 & ~n2315 ) | ( x8 & ~n2315 ) ;
  assign n2318 = n2316 & ~n2317 ;
  assign n2319 = n2313 | n2318 ;
  assign n2320 = ( n584 & ~n2308 ) | ( n584 & n2319 ) | ( ~n2308 & n2319 ) ;
  assign n2321 = ~x0 & n2320 ;
  assign n2322 = x2 & ~n2321 ;
  assign n2323 = n2307 & ~n2322 ;
  assign n2324 = x5 | n2323 ;
  assign n2325 = ( x8 & n551 ) | ( x8 & n1706 ) | ( n551 & n1706 ) ;
  assign n2326 = ( x3 & x8 ) | ( x3 & ~n2325 ) | ( x8 & ~n2325 ) ;
  assign n2327 = ( x7 & ~n551 ) | ( x7 & n2326 ) | ( ~n551 & n2326 ) ;
  assign n2328 = ( n551 & ~n2325 ) | ( n551 & n2327 ) | ( ~n2325 & n2327 ) ;
  assign n2329 = x1 & ~n2328 ;
  assign n2330 = x7 & n150 ;
  assign n2331 = x6 | n150 ;
  assign n2332 = ( x7 & x8 ) | ( x7 & n2331 ) | ( x8 & n2331 ) ;
  assign n2333 = ~n2330 & n2332 ;
  assign n2334 = x1 | n2333 ;
  assign n2335 = ( ~x1 & n2329 ) | ( ~x1 & n2334 ) | ( n2329 & n2334 ) ;
  assign n2336 = x2 & ~n2335 ;
  assign n2337 = x6 & ~n21 ;
  assign n2338 = ( x3 & ~n21 ) | ( x3 & n2337 ) | ( ~n21 & n2337 ) ;
  assign n2339 = ~x1 & n2338 ;
  assign n2340 = x2 | n2339 ;
  assign n2341 = ~n2336 & n2340 ;
  assign n2342 = ~x0 & n2341 ;
  assign n2343 = x5 & ~n2342 ;
  assign n2344 = n2324 & ~n2343 ;
  assign n2345 = ( ~x4 & n2291 ) | ( ~x4 & n2344 ) | ( n2291 & n2344 ) ;
  assign n2346 = n2292 | n2345 ;
  assign n2347 = x2 & x6 ;
  assign n2348 = ( x4 & x8 ) | ( x4 & n2347 ) | ( x8 & n2347 ) ;
  assign n2349 = x4 | n2348 ;
  assign n2350 = x4 & n2348 ;
  assign n2351 = n2349 & ~n2350 ;
  assign n2352 = x5 | n2351 ;
  assign n2353 = x8 & n470 ;
  assign n2354 = ( x8 & n689 ) | ( x8 & ~n2353 ) | ( n689 & ~n2353 ) ;
  assign n2355 = x2 | n2354 ;
  assign n2356 = x5 & n2355 ;
  assign n2357 = n2352 & ~n2356 ;
  assign n2358 = x1 & ~n2357 ;
  assign n2359 = ( x2 & x4 ) | ( x2 & ~n596 ) | ( x4 & ~n596 ) ;
  assign n2360 = ( x2 & ~x6 ) | ( x2 & n596 ) | ( ~x6 & n596 ) ;
  assign n2361 = ( x4 & ~x5 ) | ( x4 & n2360 ) | ( ~x5 & n2360 ) ;
  assign n2362 = n2359 & ~n2361 ;
  assign n2363 = ~x8 & n2362 ;
  assign n2364 = x1 | n2363 ;
  assign n2365 = ~n2358 & n2364 ;
  assign n2366 = x3 & n2365 ;
  assign n2367 = ( x4 & x5 ) | ( x4 & x8 ) | ( x5 & x8 ) ;
  assign n2368 = ( ~x6 & x8 ) | ( ~x6 & n2367 ) | ( x8 & n2367 ) ;
  assign n2369 = x8 & ~n2368 ;
  assign n2370 = n2368 | n2369 ;
  assign n2371 = ( ~x8 & n2369 ) | ( ~x8 & n2370 ) | ( n2369 & n2370 ) ;
  assign n2372 = x1 & ~n2371 ;
  assign n2373 = ~x4 & n695 ;
  assign n2374 = x1 | n2373 ;
  assign n2375 = ~n2372 & n2374 ;
  assign n2376 = ~x6 & n695 ;
  assign n2377 = x1 & n539 ;
  assign n2378 = n2376 & n2377 ;
  assign n2379 = x2 & ~n2378 ;
  assign n2380 = ( n2375 & n2378 ) | ( n2375 & ~n2379 ) | ( n2378 & ~n2379 ) ;
  assign n2381 = ( x2 & x4 ) | ( x2 & ~x8 ) | ( x4 & ~x8 ) ;
  assign n2382 = ( ~x4 & x6 ) | ( ~x4 & n2381 ) | ( x6 & n2381 ) ;
  assign n2383 = ( x2 & x6 ) | ( x2 & ~n2381 ) | ( x6 & ~n2381 ) ;
  assign n2384 = n2382 & ~n2383 ;
  assign n2385 = x1 | n2384 ;
  assign n2386 = x2 & n1384 ;
  assign n2387 = x1 & ~n2386 ;
  assign n2388 = n2385 & ~n2387 ;
  assign n2389 = n2380 | n2388 ;
  assign n2390 = ~x3 & n2389 ;
  assign n2391 = n2366 | n2390 ;
  assign n2392 = x0 & n2391 ;
  assign n2393 = ( x6 & x8 ) | ( x6 & n266 ) | ( x8 & n266 ) ;
  assign n2394 = ( x5 & ~x6 ) | ( x5 & n2393 ) | ( ~x6 & n2393 ) ;
  assign n2395 = ( x5 & x8 ) | ( x5 & ~n2393 ) | ( x8 & ~n2393 ) ;
  assign n2396 = n2394 & ~n2395 ;
  assign n2397 = ( ~x1 & x4 ) | ( ~x1 & x5 ) | ( x4 & x5 ) ;
  assign n2398 = ( ~x1 & x5 ) | ( ~x1 & x6 ) | ( x5 & x6 ) ;
  assign n2399 = n2397 & ~n2398 ;
  assign n2400 = x3 & n2399 ;
  assign n2401 = ( x0 & x2 ) | ( x0 & n2400 ) | ( x2 & n2400 ) ;
  assign n2402 = ~x0 & n2401 ;
  assign n2403 = ( ~n95 & n320 ) | ( ~n95 & n2402 ) | ( n320 & n2402 ) ;
  assign n2404 = n596 & ~n2403 ;
  assign n2405 = ( n596 & n2402 ) | ( n596 & ~n2404 ) | ( n2402 & ~n2404 ) ;
  assign n2406 = n2396 | n2405 ;
  assign n2407 = ( n2391 & ~n2392 ) | ( n2391 & n2406 ) | ( ~n2392 & n2406 ) ;
  assign n2408 = n2346 | n2407 ;
  assign n2409 = ( n2224 & ~n2225 ) | ( n2224 & n2408 ) | ( ~n2225 & n2408 ) ;
  assign n2410 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n2411 = ~x5 & n2410 ;
  assign n2412 = ( ~x4 & n2410 ) | ( ~x4 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = n101 & n2412 ;
  assign n2414 = ( x1 & x3 ) | ( x1 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n2415 = ( x0 & ~x1 ) | ( x0 & n2414 ) | ( ~x1 & n2414 ) ;
  assign n2416 = ( x1 & ~x3 ) | ( x1 & n2415 ) | ( ~x3 & n2415 ) ;
  assign n2417 = ~n2414 & n2416 ;
  assign n2418 = ( ~x0 & n2415 ) | ( ~x0 & n2417 ) | ( n2415 & n2417 ) ;
  assign n2419 = ~x0 & n936 ;
  assign n2420 = n57 & n2419 ;
  assign n2421 = ( ~n2413 & n2418 ) | ( ~n2413 & n2420 ) | ( n2418 & n2420 ) ;
  assign n2422 = x2 & ~n2420 ;
  assign n2423 = ( n2413 & n2421 ) | ( n2413 & ~n2422 ) | ( n2421 & ~n2422 ) ;
  assign n2424 = n1579 & n2423 ;
  assign n2425 = ~x7 & n105 ;
  assign n2426 = ( x4 & x6 ) | ( x4 & n2425 ) | ( x6 & n2425 ) ;
  assign n2427 = ~x4 & n2426 ;
  assign n2428 = ( ~n15 & n551 ) | ( ~n15 & n2427 ) | ( n551 & n2427 ) ;
  assign n2429 = x4 & ~n2428 ;
  assign n2430 = ( x4 & n2427 ) | ( x4 & ~n2429 ) | ( n2427 & ~n2429 ) ;
  assign n2431 = x3 & ~n2430 ;
  assign n2432 = ( x4 & ~x7 ) | ( x4 & n921 ) | ( ~x7 & n921 ) ;
  assign n2433 = ( x2 & ~x7 ) | ( x2 & n921 ) | ( ~x7 & n921 ) ;
  assign n2434 = ( n539 & n2432 ) | ( n539 & ~n2433 ) | ( n2432 & ~n2433 ) ;
  assign n2435 = x6 & n2434 ;
  assign n2436 = x3 | n2435 ;
  assign n2437 = ~n2431 & n2436 ;
  assign n2438 = x8 & n2437 ;
  assign n2439 = ~n66 & n68 ;
  assign n2440 = ( x1 & ~n445 ) | ( x1 & n2439 ) | ( ~n445 & n2439 ) ;
  assign n2441 = ~x1 & n2440 ;
  assign n2442 = ( x6 & x7 ) | ( x6 & n37 ) | ( x7 & n37 ) ;
  assign n2443 = n1946 & ~n2442 ;
  assign n2444 = x1 & n2443 ;
  assign n2445 = ( ~x5 & x6 ) | ( ~x5 & n2184 ) | ( x6 & n2184 ) ;
  assign n2446 = ( ~x5 & x7 ) | ( ~x5 & n2184 ) | ( x7 & n2184 ) ;
  assign n2447 = ( n551 & n2445 ) | ( n551 & ~n2446 ) | ( n2445 & ~n2446 ) ;
  assign n2448 = x1 | n2447 ;
  assign n2449 = ( ~x1 & n2444 ) | ( ~x1 & n2448 ) | ( n2444 & n2448 ) ;
  assign n2450 = x8 & ~n2449 ;
  assign n2451 = ( ~x3 & n572 ) | ( ~x3 & n1874 ) | ( n572 & n1874 ) ;
  assign n2452 = ( x6 & n1874 ) | ( x6 & ~n2451 ) | ( n1874 & ~n2451 ) ;
  assign n2453 = ( x3 & n2451 ) | ( x3 & ~n2452 ) | ( n2451 & ~n2452 ) ;
  assign n2454 = x5 & n2453 ;
  assign n2455 = x8 | n2454 ;
  assign n2456 = ~n2450 & n2455 ;
  assign n2457 = x2 & n2456 ;
  assign n2458 = ( x3 & n584 ) | ( x3 & n1856 ) | ( n584 & n1856 ) ;
  assign n2459 = ~x3 & n2458 ;
  assign n2460 = ( x1 & x7 ) | ( x1 & n898 ) | ( x7 & n898 ) ;
  assign n2461 = ( x6 & x7 ) | ( x6 & ~n2460 ) | ( x7 & ~n2460 ) ;
  assign n2462 = x5 & n2461 ;
  assign n2463 = ( x1 & ~n2460 ) | ( x1 & n2462 ) | ( ~n2460 & n2462 ) ;
  assign n2464 = ( x3 & n2459 ) | ( x3 & n2463 ) | ( n2459 & n2463 ) ;
  assign n2465 = x8 & ~n2464 ;
  assign n2466 = ( x8 & n2459 ) | ( x8 & ~n2465 ) | ( n2459 & ~n2465 ) ;
  assign n2467 = ( x1 & ~x3 ) | ( x1 & x8 ) | ( ~x3 & x8 ) ;
  assign n2468 = ( x1 & ~x7 ) | ( x1 & n2467 ) | ( ~x7 & n2467 ) ;
  assign n2469 = x1 & ~n2468 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = ( ~x1 & n2469 ) | ( ~x1 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = ( x5 & x6 ) | ( x5 & n2471 ) | ( x6 & n2471 ) ;
  assign n2473 = ( ~n596 & n2466 ) | ( ~n596 & n2472 ) | ( n2466 & n2472 ) ;
  assign n2474 = x2 | n2473 ;
  assign n2475 = ( ~x2 & n2457 ) | ( ~x2 & n2474 ) | ( n2457 & n2474 ) ;
  assign n2476 = x4 & n2475 ;
  assign n2477 = ( x2 & ~x5 ) | ( x2 & n2414 ) | ( ~x5 & n2414 ) ;
  assign n2478 = x5 & n2477 ;
  assign n2479 = n2477 & ~n2478 ;
  assign n2480 = ( x5 & ~n2478 ) | ( x5 & n2479 ) | ( ~n2478 & n2479 ) ;
  assign n2481 = n584 & ~n2480 ;
  assign n2482 = ( n575 & ~n2480 ) | ( n575 & n2481 ) | ( ~n2480 & n2481 ) ;
  assign n2483 = ( x1 & x8 ) | ( x1 & ~n2237 ) | ( x8 & ~n2237 ) ;
  assign n2484 = ( ~x5 & x6 ) | ( ~x5 & n2483 ) | ( x6 & n2483 ) ;
  assign n2485 = n2237 & n2484 ;
  assign n2486 = ( ~n2483 & n2484 ) | ( ~n2483 & n2485 ) | ( n2484 & n2485 ) ;
  assign n2487 = ~x1 & n584 ;
  assign n2488 = ~x5 & n2487 ;
  assign n2489 = x7 & ~n2488 ;
  assign n2490 = ( n2486 & n2488 ) | ( n2486 & ~n2489 ) | ( n2488 & ~n2489 ) ;
  assign n2491 = x3 & ~n2490 ;
  assign n2492 = x1 & n553 ;
  assign n2493 = x3 | n2492 ;
  assign n2494 = ~n2491 & n2493 ;
  assign n2495 = ~x2 & n2494 ;
  assign n2496 = ( x8 & n74 ) | ( x8 & ~n811 ) | ( n74 & ~n811 ) ;
  assign n2497 = ( ~x6 & x7 ) | ( ~x6 & n213 ) | ( x7 & n213 ) ;
  assign n2498 = ( ~x3 & x6 ) | ( ~x3 & n213 ) | ( x6 & n213 ) ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = x1 & ~n2499 ;
  assign n2501 = x8 & n2500 ;
  assign n2502 = ( n811 & n2496 ) | ( n811 & n2501 ) | ( n2496 & n2501 ) ;
  assign n2503 = x1 & n584 ;
  assign n2504 = n37 & n2503 ;
  assign n2505 = n2502 | n2504 ;
  assign n2506 = x2 & n2505 ;
  assign n2507 = n2495 | n2506 ;
  assign n2508 = n2482 | n2507 ;
  assign n2509 = ~x4 & n2508 ;
  assign n2510 = n2476 | n2509 ;
  assign n2511 = n2441 | n2510 ;
  assign n2512 = ( n2437 & ~n2438 ) | ( n2437 & n2511 ) | ( ~n2438 & n2511 ) ;
  assign n2513 = x0 & n2512 ;
  assign n2514 = n1638 & ~n1984 ;
  assign n2515 = n1259 & n2514 ;
  assign n2516 = x4 & n66 ;
  assign n2517 = ( n1305 & n1350 ) | ( n1305 & ~n2516 ) | ( n1350 & ~n2516 ) ;
  assign n2518 = ( ~x8 & n2515 ) | ( ~x8 & n2517 ) | ( n2515 & n2517 ) ;
  assign n2519 = x7 & ~n2518 ;
  assign n2520 = ( x7 & n2515 ) | ( x7 & ~n2519 ) | ( n2515 & ~n2519 ) ;
  assign n2521 = x5 & n2520 ;
  assign n2522 = ( x4 & n145 ) | ( x4 & n672 ) | ( n145 & n672 ) ;
  assign n2523 = ~x4 & n2522 ;
  assign n2524 = n2521 | n2523 ;
  assign n2525 = ( ~x0 & n2521 ) | ( ~x0 & n2524 ) | ( n2521 & n2524 ) ;
  assign n2526 = x1 | n2525 ;
  assign n2527 = ( x3 & x4 ) | ( x3 & n306 ) | ( x4 & n306 ) ;
  assign n2528 = ( ~x2 & x4 ) | ( ~x2 & n306 ) | ( x4 & n306 ) ;
  assign n2529 = ( n66 & ~n2527 ) | ( n66 & n2528 ) | ( ~n2527 & n2528 ) ;
  assign n2530 = ~x8 & n22 ;
  assign n2531 = n842 & n2530 ;
  assign n2532 = x5 & ~n2531 ;
  assign n2533 = ( n2529 & ~n2531 ) | ( n2529 & n2532 ) | ( ~n2531 & n2532 ) ;
  assign n2534 = n27 & n284 ;
  assign n2535 = x7 | n2534 ;
  assign n2536 = ( ~n2533 & n2534 ) | ( ~n2533 & n2535 ) | ( n2534 & n2535 ) ;
  assign n2537 = ~x0 & n2536 ;
  assign n2538 = x1 & ~n2537 ;
  assign n2539 = n2526 & ~n2538 ;
  assign n2540 = n885 | n2539 ;
  assign n2541 = ( n2512 & ~n2513 ) | ( n2512 & n2540 ) | ( ~n2513 & n2540 ) ;
  assign n2542 = ( x0 & ~x3 ) | ( x0 & n2530 ) | ( ~x3 & n2530 ) ;
  assign n2543 = ( x4 & ~x8 ) | ( x4 & n636 ) | ( ~x8 & n636 ) ;
  assign n2544 = x4 & ~n2543 ;
  assign n2545 = n2543 | n2544 ;
  assign n2546 = ( ~x4 & n2544 ) | ( ~x4 & n2545 ) | ( n2544 & n2545 ) ;
  assign n2547 = ( x0 & x3 ) | ( x0 & ~n2546 ) | ( x3 & ~n2546 ) ;
  assign n2548 = n2542 & ~n2547 ;
  assign n2549 = x5 & n729 ;
  assign n2550 = ( x0 & n192 ) | ( x0 & n2549 ) | ( n192 & n2549 ) ;
  assign n2551 = ~x0 & n2550 ;
  assign n2552 = ~x5 & n1537 ;
  assign n2553 = ( n1537 & ~n1872 ) | ( n1537 & n2552 ) | ( ~n1872 & n2552 ) ;
  assign n2554 = ( x1 & n1350 ) | ( x1 & n2553 ) | ( n1350 & n2553 ) ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = ( ~n2548 & n2551 ) | ( ~n2548 & n2555 ) | ( n2551 & n2555 ) ;
  assign n2557 = x1 & ~n2555 ;
  assign n2558 = ( n2548 & n2556 ) | ( n2548 & ~n2557 ) | ( n2556 & ~n2557 ) ;
  assign n2559 = x2 | n2558 ;
  assign n2560 = ( x3 & x5 ) | ( x3 & ~x8 ) | ( x5 & ~x8 ) ;
  assign n2561 = ( ~x3 & x6 ) | ( ~x3 & n2560 ) | ( x6 & n2560 ) ;
  assign n2562 = ( x5 & x6 ) | ( x5 & ~n2560 ) | ( x6 & ~n2560 ) ;
  assign n2563 = n2561 & ~n2562 ;
  assign n2564 = ( x1 & ~x4 ) | ( x1 & n2563 ) | ( ~x4 & n2563 ) ;
  assign n2565 = ( x3 & x5 ) | ( x3 & x8 ) | ( x5 & x8 ) ;
  assign n2566 = ( x3 & x6 ) | ( x3 & ~n2565 ) | ( x6 & ~n2565 ) ;
  assign n2567 = ( ~x5 & x6 ) | ( ~x5 & n2565 ) | ( x6 & n2565 ) ;
  assign n2568 = ~n2566 & n2567 ;
  assign n2569 = ( x1 & x4 ) | ( x1 & ~n2568 ) | ( x4 & ~n2568 ) ;
  assign n2570 = n2564 & ~n2569 ;
  assign n2571 = ( ~x1 & n26 ) | ( ~x1 & n2570 ) | ( n26 & n2570 ) ;
  assign n2572 = n983 | n2571 ;
  assign n2573 = ( ~n983 & n2570 ) | ( ~n983 & n2572 ) | ( n2570 & n2572 ) ;
  assign n2574 = ~x0 & n2573 ;
  assign n2575 = x2 & ~n2574 ;
  assign n2576 = n2559 & ~n2575 ;
  assign n2577 = n2541 | n2576 ;
  assign n2578 = ( n2423 & ~n2424 ) | ( n2423 & n2577 ) | ( ~n2424 & n2577 ) ;
  assign n2579 = ( x5 & ~x8 ) | ( x5 & n1618 ) | ( ~x8 & n1618 ) ;
  assign n2580 = ( x1 & x4 ) | ( x1 & n2579 ) | ( x4 & n2579 ) ;
  assign n2581 = ~n1618 & n2580 ;
  assign n2582 = ( ~n2579 & n2580 ) | ( ~n2579 & n2581 ) | ( n2580 & n2581 ) ;
  assign n2583 = x3 & ~n2582 ;
  assign n2584 = ~x1 & n1536 ;
  assign n2585 = x3 | n2584 ;
  assign n2586 = ~n2583 & n2585 ;
  assign n2587 = ( ~x0 & x2 ) | ( ~x0 & n2586 ) | ( x2 & n2586 ) ;
  assign n2588 = x3 & ~n1633 ;
  assign n2589 = ~x5 & n2588 ;
  assign n2590 = ( x8 & ~n1633 ) | ( x8 & n2588 ) | ( ~n1633 & n2588 ) ;
  assign n2591 = ( x1 & n2589 ) | ( x1 & n2590 ) | ( n2589 & n2590 ) ;
  assign n2592 = x4 | n2591 ;
  assign n2593 = x8 | n1387 ;
  assign n2594 = x1 & ~n2593 ;
  assign n2595 = x4 & ~n2594 ;
  assign n2596 = n2592 & ~n2595 ;
  assign n2597 = ( x0 & x2 ) | ( x0 & ~n2596 ) | ( x2 & ~n2596 ) ;
  assign n2598 = n2587 & ~n2597 ;
  assign n2599 = ( x5 & ~n320 ) | ( x5 & n458 ) | ( ~n320 & n458 ) ;
  assign n2600 = n320 & n2599 ;
  assign n2601 = n2598 | n2600 ;
  assign n2602 = ( ~x6 & x7 ) | ( ~x6 & n2601 ) | ( x7 & n2601 ) ;
  assign n2603 = ( n551 & n2601 ) | ( n551 & ~n2602 ) | ( n2601 & ~n2602 ) ;
  assign n2604 = ( ~x6 & x8 ) | ( ~x6 & n218 ) | ( x8 & n218 ) ;
  assign n2605 = x8 & ~n2604 ;
  assign n2606 = n2604 | n2605 ;
  assign n2607 = ( ~x8 & n2605 ) | ( ~x8 & n2606 ) | ( n2605 & n2606 ) ;
  assign n2608 = x4 & n2607 ;
  assign n2609 = x1 & ~n2608 ;
  assign n2610 = ~n58 & n60 ;
  assign n2611 = x1 | n2610 ;
  assign n2612 = ~n2609 & n2611 ;
  assign n2613 = ( ~x0 & x2 ) | ( ~x0 & n2612 ) | ( x2 & n2612 ) ;
  assign n2614 = ( x6 & ~x7 ) | ( x6 & n998 ) | ( ~x7 & n998 ) ;
  assign n2615 = x6 & ~n2614 ;
  assign n2616 = n2614 | n2615 ;
  assign n2617 = ( ~x6 & n2615 ) | ( ~x6 & n2616 ) | ( n2615 & n2616 ) ;
  assign n2618 = x1 | n2617 ;
  assign n2619 = x1 & ~n1171 ;
  assign n2620 = n2618 & ~n2619 ;
  assign n2621 = x3 | n2620 ;
  assign n2622 = ( ~x4 & x7 ) | ( ~x4 & n1489 ) | ( x7 & n1489 ) ;
  assign n2623 = ( ~x7 & x8 ) | ( ~x7 & n1489 ) | ( x8 & n1489 ) ;
  assign n2624 = n2622 & n2623 ;
  assign n2625 = x1 & n2624 ;
  assign n2626 = x3 & ~n2625 ;
  assign n2627 = n2621 & ~n2626 ;
  assign n2628 = ( x0 & x2 ) | ( x0 & ~n2627 ) | ( x2 & ~n2627 ) ;
  assign n2629 = n2613 & ~n2628 ;
  assign n2630 = ( n10 & n99 ) | ( n10 & n2629 ) | ( n99 & n2629 ) ;
  assign n2631 = n445 | n2630 ;
  assign n2632 = ( ~n445 & n2629 ) | ( ~n445 & n2631 ) | ( n2629 & n2631 ) ;
  assign n2633 = ( x0 & x3 ) | ( x0 & ~x4 ) | ( x3 & ~x4 ) ;
  assign n2634 = ( x0 & x3 ) | ( x0 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n2635 = n2633 & n2634 ;
  assign n2636 = x5 | n2635 ;
  assign n2637 = ( ~n2633 & n2635 ) | ( ~n2633 & n2636 ) | ( n2635 & n2636 ) ;
  assign n2638 = ( ~x2 & x6 ) | ( ~x2 & n2637 ) | ( x6 & n2637 ) ;
  assign n2639 = ( x2 & n1263 ) | ( x2 & n1387 ) | ( n1263 & n1387 ) ;
  assign n2640 = ~n1387 & n2639 ;
  assign n2641 = x6 & n2640 ;
  assign n2642 = ( ~n2637 & n2638 ) | ( ~n2637 & n2641 ) | ( n2638 & n2641 ) ;
  assign n2643 = ~x3 & n2191 ;
  assign n2644 = ( x2 & x5 ) | ( x2 & ~n2643 ) | ( x5 & ~n2643 ) ;
  assign n2645 = ( n2191 & n2643 ) | ( n2191 & ~n2644 ) | ( n2643 & ~n2644 ) ;
  assign n2646 = ( ~x0 & n2642 ) | ( ~x0 & n2645 ) | ( n2642 & n2645 ) ;
  assign n2647 = x4 & ~n2646 ;
  assign n2648 = ( x4 & n2642 ) | ( x4 & ~n2647 ) | ( n2642 & ~n2647 ) ;
  assign n2649 = ( x2 & x5 ) | ( x2 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n2650 = ~n232 & n2649 ;
  assign n2651 = ~x4 & n2650 ;
  assign n2652 = ( x0 & ~x6 ) | ( x0 & n2651 ) | ( ~x6 & n2651 ) ;
  assign n2653 = ~x0 & n2652 ;
  assign n2654 = x7 | n2653 ;
  assign n2655 = ( n2648 & n2653 ) | ( n2648 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = x1 | n2655 ;
  assign n2657 = ( x4 & x5 ) | ( x4 & x7 ) | ( x5 & x7 ) ;
  assign n2658 = n1984 & ~n2657 ;
  assign n2659 = ( x2 & ~x6 ) | ( x2 & n2658 ) | ( ~x6 & n2658 ) ;
  assign n2660 = x4 & n36 ;
  assign n2661 = n130 & n2660 ;
  assign n2662 = ~x6 & n2661 ;
  assign n2663 = ( ~x2 & n2659 ) | ( ~x2 & n2662 ) | ( n2659 & n2662 ) ;
  assign n2664 = ~x0 & n2663 ;
  assign n2665 = x1 & ~n2664 ;
  assign n2666 = n2656 & ~n2665 ;
  assign n2667 = ( ~x3 & x5 ) | ( ~x3 & n1629 ) | ( x5 & n1629 ) ;
  assign n2668 = ( x1 & x7 ) | ( x1 & n2667 ) | ( x7 & n2667 ) ;
  assign n2669 = ~n1629 & n2668 ;
  assign n2670 = ( ~n2667 & n2668 ) | ( ~n2667 & n2669 ) | ( n2668 & n2669 ) ;
  assign n2671 = x4 & n2670 ;
  assign n2672 = ~x0 & n2671 ;
  assign n2673 = ( ~x4 & n130 ) | ( ~x4 & n2672 ) | ( n130 & n2672 ) ;
  assign n2674 = n1357 & ~n2673 ;
  assign n2675 = ( n1357 & n2672 ) | ( n1357 & ~n2674 ) | ( n2672 & ~n2674 ) ;
  assign n2676 = ~n357 & n789 ;
  assign n2677 = ( x5 & ~n101 ) | ( x5 & n1706 ) | ( ~n101 & n1706 ) ;
  assign n2678 = n101 & n2677 ;
  assign n2679 = ( x3 & ~x5 ) | ( x3 & x7 ) | ( ~x5 & x7 ) ;
  assign n2680 = ( x1 & x5 ) | ( x1 & n2679 ) | ( x5 & n2679 ) ;
  assign n2681 = ( x5 & x7 ) | ( x5 & ~n2680 ) | ( x7 & ~n2680 ) ;
  assign n2682 = n2679 | n2681 ;
  assign n2683 = ( x1 & ~n2680 ) | ( x1 & n2682 ) | ( ~n2680 & n2682 ) ;
  assign n2684 = ( x0 & ~x4 ) | ( x0 & n2683 ) | ( ~x4 & n2683 ) ;
  assign n2685 = ( x3 & ~x5 ) | ( x3 & n1629 ) | ( ~x5 & n1629 ) ;
  assign n2686 = x3 & ~n2685 ;
  assign n2687 = n2685 | n2686 ;
  assign n2688 = ( ~x3 & n2686 ) | ( ~x3 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = ( x0 & x4 ) | ( x0 & ~n2688 ) | ( x4 & ~n2688 ) ;
  assign n2690 = n2684 | n2689 ;
  assign n2691 = ~n2678 & n2690 ;
  assign n2692 = ~n2676 & n2691 ;
  assign n2693 = ~x6 & n2692 ;
  assign n2694 = ( x1 & x5 ) | ( x1 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n2695 = ( ~x1 & x7 ) | ( ~x1 & n2694 ) | ( x7 & n2694 ) ;
  assign n2696 = ( ~x3 & x7 ) | ( ~x3 & n2695 ) | ( x7 & n2695 ) ;
  assign n2697 = ( ~n37 & n2694 ) | ( ~n37 & n2696 ) | ( n2694 & n2696 ) ;
  assign n2698 = ~x4 & n2697 ;
  assign n2699 = n74 & n130 ;
  assign n2700 = x4 & ~n2699 ;
  assign n2701 = n2698 | n2700 ;
  assign n2702 = x0 | n2701 ;
  assign n2703 = x6 & n2702 ;
  assign n2704 = n2693 | n2703 ;
  assign n2705 = x8 & n2704 ;
  assign n2706 = ( ~x3 & x5 ) | ( ~x3 & n394 ) | ( x5 & n394 ) ;
  assign n2707 = ( x4 & x5 ) | ( x4 & ~n394 ) | ( x5 & ~n394 ) ;
  assign n2708 = ( ~x3 & x7 ) | ( ~x3 & n2707 ) | ( x7 & n2707 ) ;
  assign n2709 = ~n2706 & n2708 ;
  assign n2710 = x1 & n2709 ;
  assign n2711 = ( x3 & x5 ) | ( x3 & ~n1563 ) | ( x5 & ~n1563 ) ;
  assign n2712 = ( x4 & ~x7 ) | ( x4 & n2711 ) | ( ~x7 & n2711 ) ;
  assign n2713 = n1563 & n2712 ;
  assign n2714 = ( ~n2711 & n2712 ) | ( ~n2711 & n2713 ) | ( n2712 & n2713 ) ;
  assign n2715 = x1 | n2714 ;
  assign n2716 = ( ~x1 & n2710 ) | ( ~x1 & n2715 ) | ( n2710 & n2715 ) ;
  assign n2717 = x6 & ~n2716 ;
  assign n2718 = x7 & ~n26 ;
  assign n2719 = ( ~n738 & n764 ) | ( ~n738 & n2718 ) | ( n764 & n2718 ) ;
  assign n2720 = x1 & ~n2719 ;
  assign n2721 = x6 | n2720 ;
  assign n2722 = ~n2717 & n2721 ;
  assign n2723 = ~x0 & n2722 ;
  assign n2724 = x8 | n2723 ;
  assign n2725 = ~n2705 & n2724 ;
  assign n2726 = n762 & ~n2725 ;
  assign n2727 = ( n2675 & n2725 ) | ( n2675 & ~n2726 ) | ( n2725 & ~n2726 ) ;
  assign n2728 = x2 | n2727 ;
  assign n2729 = n59 | n68 ;
  assign n2730 = ( n52 & n59 ) | ( n52 & n2729 ) | ( n59 & n2729 ) ;
  assign n2731 = x1 & ~n2730 ;
  assign n2732 = x5 & n575 ;
  assign n2733 = x1 | n2732 ;
  assign n2734 = ~n2731 & n2733 ;
  assign n2735 = ( x3 & ~x6 ) | ( x3 & x8 ) | ( ~x6 & x8 ) ;
  assign n2736 = ( ~x3 & x6 ) | ( ~x3 & n2735 ) | ( x6 & n2735 ) ;
  assign n2737 = ~x1 & n2735 ;
  assign n2738 = ( ~x8 & n2735 ) | ( ~x8 & n2737 ) | ( n2735 & n2737 ) ;
  assign n2739 = n2736 | n2738 ;
  assign n2740 = ( x5 & n2734 ) | ( x5 & ~n2739 ) | ( n2734 & ~n2739 ) ;
  assign n2741 = x7 & ~n2740 ;
  assign n2742 = ( x7 & n2734 ) | ( x7 & ~n2741 ) | ( n2734 & ~n2741 ) ;
  assign n2743 = ~x4 & n2742 ;
  assign n2744 = ( x1 & x5 ) | ( x1 & ~n68 ) | ( x5 & ~n68 ) ;
  assign n2745 = ( ~x1 & x7 ) | ( ~x1 & n2744 ) | ( x7 & n2744 ) ;
  assign n2746 = ( ~x5 & x8 ) | ( ~x5 & n2745 ) | ( x8 & n2745 ) ;
  assign n2747 = n2744 & n2746 ;
  assign n2748 = ( ~x3 & x6 ) | ( ~x3 & n2747 ) | ( x6 & n2747 ) ;
  assign n2749 = ( x1 & x7 ) | ( x1 & n614 ) | ( x7 & n614 ) ;
  assign n2750 = ( x3 & ~x7 ) | ( x3 & n2749 ) | ( ~x7 & n2749 ) ;
  assign n2751 = ( x1 & x3 ) | ( x1 & ~n2749 ) | ( x3 & ~n2749 ) ;
  assign n2752 = n2750 & ~n2751 ;
  assign n2753 = ~x6 & n2752 ;
  assign n2754 = ( n2747 & ~n2748 ) | ( n2747 & n2753 ) | ( ~n2748 & n2753 ) ;
  assign n2755 = ( x1 & x7 ) | ( x1 & x8 ) | ( x7 & x8 ) ;
  assign n2756 = ( ~x3 & x8 ) | ( ~x3 & n2755 ) | ( x8 & n2755 ) ;
  assign n2757 = x8 & ~n2756 ;
  assign n2758 = n2756 | n2757 ;
  assign n2759 = ( ~x8 & n2757 ) | ( ~x8 & n2758 ) | ( n2757 & n2758 ) ;
  assign n2760 = ( x5 & x6 ) | ( x5 & ~n2759 ) | ( x6 & ~n2759 ) ;
  assign n2761 = ( x1 & x7 ) | ( x1 & ~n1528 ) | ( x7 & ~n1528 ) ;
  assign n2762 = x1 & ~n2761 ;
  assign n2763 = ( x7 & ~n2761 ) | ( x7 & n2762 ) | ( ~n2761 & n2762 ) ;
  assign n2764 = x6 & n2763 ;
  assign n2765 = ( n2759 & n2760 ) | ( n2759 & n2764 ) | ( n2760 & n2764 ) ;
  assign n2766 = n2754 | n2765 ;
  assign n2767 = x4 & n2766 ;
  assign n2768 = n2743 | n2767 ;
  assign n2769 = ~x0 & n2768 ;
  assign n2770 = x2 & ~n2769 ;
  assign n2771 = n2728 & ~n2770 ;
  assign n2772 = n2666 | n2771 ;
  assign n2773 = ( ~n2603 & n2632 ) | ( ~n2603 & n2772 ) | ( n2632 & n2772 ) ;
  assign n2774 = n2603 | n2773 ;
  assign n2775 = ~x3 & n447 ;
  assign n2776 = n98 & ~n2775 ;
  assign n2777 = x2 & n101 ;
  assign n2778 = ( x3 & x8 ) | ( x3 & n2777 ) | ( x8 & n2777 ) ;
  assign n2779 = ~x8 & n2778 ;
  assign n2780 = ( x2 & x8 ) | ( x2 & ~n1484 ) | ( x8 & ~n1484 ) ;
  assign n2781 = ( x2 & x5 ) | ( x2 & ~n1484 ) | ( x5 & ~n1484 ) ;
  assign n2782 = ( n613 & n2780 ) | ( n613 & ~n2781 ) | ( n2780 & ~n2781 ) ;
  assign n2783 = ( ~x0 & x3 ) | ( ~x0 & n2782 ) | ( x3 & n2782 ) ;
  assign n2784 = ( x1 & ~x5 ) | ( x1 & x8 ) | ( ~x5 & x8 ) ;
  assign n2785 = ~x1 & n2784 ;
  assign n2786 = ( x2 & x8 ) | ( x2 & ~n2785 ) | ( x8 & ~n2785 ) ;
  assign n2787 = ( n2784 & n2785 ) | ( n2784 & ~n2786 ) | ( n2785 & ~n2786 ) ;
  assign n2788 = ( x0 & x3 ) | ( x0 & ~n2787 ) | ( x3 & ~n2787 ) ;
  assign n2789 = n2783 & ~n2788 ;
  assign n2790 = n2779 | n2789 ;
  assign n2791 = ( n98 & ~n2776 ) | ( n98 & n2790 ) | ( ~n2776 & n2790 ) ;
  assign n2792 = x4 & n2791 ;
  assign n2793 = ( x0 & x5 ) | ( x0 & x8 ) | ( x5 & x8 ) ;
  assign n2794 = ( ~x0 & x3 ) | ( ~x0 & n2793 ) | ( x3 & n2793 ) ;
  assign n2795 = ( x5 & x8 ) | ( x5 & n2794 ) | ( x8 & n2794 ) ;
  assign n2796 = n2793 & ~n2795 ;
  assign n2797 = ( n2794 & ~n2795 ) | ( n2794 & n2796 ) | ( ~n2795 & n2796 ) ;
  assign n2798 = ( x1 & x2 ) | ( x1 & n2797 ) | ( x2 & n2797 ) ;
  assign n2799 = n101 & ~n2593 ;
  assign n2800 = ~x2 & n2799 ;
  assign n2801 = ( n2797 & ~n2798 ) | ( n2797 & n2800 ) | ( ~n2798 & n2800 ) ;
  assign n2802 = ( x5 & ~n106 ) | ( x5 & n1530 ) | ( ~n106 & n1530 ) ;
  assign n2803 = n106 & n2802 ;
  assign n2804 = n2801 | n2803 ;
  assign n2805 = ~x4 & n2804 ;
  assign n2806 = n2792 | n2805 ;
  assign n2807 = ( x6 & x7 ) | ( x6 & ~n2806 ) | ( x7 & ~n2806 ) ;
  assign n2808 = x6 & ~n2807 ;
  assign n2809 = ( x7 & ~n2807 ) | ( x7 & n2808 ) | ( ~n2807 & n2808 ) ;
  assign n2810 = x0 & ~x7 ;
  assign n2811 = x4 & ~n2810 ;
  assign n2812 = ( n68 & n689 ) | ( n68 & ~n2811 ) | ( n689 & ~n2811 ) ;
  assign n2813 = x6 & ~n2812 ;
  assign n2814 = x0 | n880 ;
  assign n2815 = ~x6 & n2814 ;
  assign n2816 = n2813 | n2815 ;
  assign n2817 = ~x3 & n2816 ;
  assign n2818 = ~x8 & n242 ;
  assign n2819 = ( x6 & x8 ) | ( x6 & ~n242 ) | ( x8 & ~n242 ) ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = ( x8 & n2818 ) | ( x8 & n2820 ) | ( n2818 & n2820 ) ;
  assign n2822 = x0 | n2821 ;
  assign n2823 = x3 & n2822 ;
  assign n2824 = n2817 | n2823 ;
  assign n2825 = ~x2 & n2824 ;
  assign n2826 = ( ~x7 & x8 ) | ( ~x7 & n1575 ) | ( x8 & n1575 ) ;
  assign n2827 = ( ~x4 & x8 ) | ( ~x4 & n1575 ) | ( x8 & n1575 ) ;
  assign n2828 = ( n83 & ~n2826 ) | ( n83 & n2827 ) | ( ~n2826 & n2827 ) ;
  assign n2829 = x6 | n2828 ;
  assign n2830 = ~x4 & n21 ;
  assign n2831 = x6 & ~n2830 ;
  assign n2832 = n2829 & ~n2831 ;
  assign n2833 = ~x0 & n2832 ;
  assign n2834 = x2 & ~n2833 ;
  assign n2835 = n2825 | n2834 ;
  assign n2836 = ~x1 & n2835 ;
  assign n2837 = ( x3 & x6 ) | ( x3 & x7 ) | ( x6 & x7 ) ;
  assign n2838 = ( x3 & x8 ) | ( x3 & ~n2837 ) | ( x8 & ~n2837 ) ;
  assign n2839 = ( ~x3 & x6 ) | ( ~x3 & n2838 ) | ( x6 & n2838 ) ;
  assign n2840 = n2837 | n2839 ;
  assign n2841 = ( ~x8 & n2838 ) | ( ~x8 & n2840 ) | ( n2838 & n2840 ) ;
  assign n2842 = x4 & ~n2841 ;
  assign n2843 = ( x3 & ~n451 ) | ( x3 & n1656 ) | ( ~n451 & n1656 ) ;
  assign n2844 = x4 | n2843 ;
  assign n2845 = ( ~x4 & n2842 ) | ( ~x4 & n2844 ) | ( n2842 & n2844 ) ;
  assign n2846 = x2 & n2845 ;
  assign n2847 = x8 & ~n145 ;
  assign n2848 = ~x6 & n2847 ;
  assign n2849 = ( x3 & ~n145 ) | ( x3 & n2847 ) | ( ~n145 & n2847 ) ;
  assign n2850 = ( ~x7 & n2848 ) | ( ~x7 & n2849 ) | ( n2848 & n2849 ) ;
  assign n2851 = x4 & ~n2850 ;
  assign n2852 = ( x3 & x7 ) | ( x3 & n762 ) | ( x7 & n762 ) ;
  assign n2853 = x3 & ~n2852 ;
  assign n2854 = ( x7 & ~n2852 ) | ( x7 & n2853 ) | ( ~n2852 & n2853 ) ;
  assign n2855 = ~x4 & n2854 ;
  assign n2856 = ( x4 & ~n2851 ) | ( x4 & n2855 ) | ( ~n2851 & n2855 ) ;
  assign n2857 = x2 | n2856 ;
  assign n2858 = ( ~x2 & n2846 ) | ( ~x2 & n2857 ) | ( n2846 & n2857 ) ;
  assign n2859 = ~x0 & n2858 ;
  assign n2860 = x1 & ~n2859 ;
  assign n2861 = n2836 | n2860 ;
  assign n2862 = x5 & n2861 ;
  assign n2863 = ( ~x1 & x3 ) | ( ~x1 & x6 ) | ( x3 & x6 ) ;
  assign n2864 = x1 & n2863 ;
  assign n2865 = ( ~n1420 & n2863 ) | ( ~n1420 & n2864 ) | ( n2863 & n2864 ) ;
  assign n2866 = x3 | x6 ;
  assign n2867 = ( ~x3 & x7 ) | ( ~x3 & n2866 ) | ( x7 & n2866 ) ;
  assign n2868 = ( x7 & x8 ) | ( x7 & n2866 ) | ( x8 & n2866 ) ;
  assign n2869 = ( n2309 & n2867 ) | ( n2309 & ~n2868 ) | ( n2867 & ~n2868 ) ;
  assign n2870 = x2 & n2869 ;
  assign n2871 = x3 & n258 ;
  assign n2872 = x2 | n2871 ;
  assign n2873 = ~n2870 & n2872 ;
  assign n2874 = x1 & ~n2873 ;
  assign n2875 = x7 & ~n842 ;
  assign n2876 = ( ~n572 & n2866 ) | ( ~n572 & n2875 ) | ( n2866 & n2875 ) ;
  assign n2877 = x8 | n2876 ;
  assign n2878 = ~x1 & n2877 ;
  assign n2879 = n2874 | n2878 ;
  assign n2880 = ( n10 & n447 ) | ( n10 & ~n1803 ) | ( n447 & ~n1803 ) ;
  assign n2881 = n2879 & ~n2880 ;
  assign n2882 = ( ~n2865 & n2879 ) | ( ~n2865 & n2881 ) | ( n2879 & n2881 ) ;
  assign n2883 = x4 & ~n2882 ;
  assign n2884 = ( ~x6 & x8 ) | ( ~x6 & n1784 ) | ( x8 & n1784 ) ;
  assign n2885 = x8 & ~n2884 ;
  assign n2886 = n2884 | n2885 ;
  assign n2887 = ( ~x8 & n2885 ) | ( ~x8 & n2886 ) | ( n2885 & n2886 ) ;
  assign n2888 = ( ~x1 & x3 ) | ( ~x1 & n2887 ) | ( x3 & n2887 ) ;
  assign n2889 = ( n145 & n715 ) | ( n145 & ~n2347 ) | ( n715 & ~n2347 ) ;
  assign n2890 = ( x7 & n145 ) | ( x7 & n2889 ) | ( n145 & n2889 ) ;
  assign n2891 = ( x1 & x3 ) | ( x1 & n2890 ) | ( x3 & n2890 ) ;
  assign n2892 = n2888 & n2891 ;
  assign n2893 = x3 | n451 ;
  assign n2894 = ( x1 & x2 ) | ( x1 & ~n2893 ) | ( x2 & ~n2893 ) ;
  assign n2895 = ~x1 & n2894 ;
  assign n2896 = n2892 | n2895 ;
  assign n2897 = ~x4 & n2896 ;
  assign n2898 = n2883 | n2897 ;
  assign n2899 = ~x0 & n2898 ;
  assign n2900 = x5 | n2899 ;
  assign n2901 = ~n2862 & n2900 ;
  assign n2902 = ( x0 & x4 ) | ( x0 & n171 ) | ( x4 & n171 ) ;
  assign n2903 = ( x4 & x7 ) | ( x4 & ~n2902 ) | ( x7 & ~n2902 ) ;
  assign n2904 = ( x0 & ~x5 ) | ( x0 & n2903 ) | ( ~x5 & n2903 ) ;
  assign n2905 = ~n2902 & n2904 ;
  assign n2906 = x1 | n2905 ;
  assign n2907 = ~x0 & n405 ;
  assign n2908 = x1 & ~n2907 ;
  assign n2909 = n2906 & ~n2908 ;
  assign n2910 = x2 | n2909 ;
  assign n2911 = ( ~x1 & x4 ) | ( ~x1 & n1033 ) | ( x4 & n1033 ) ;
  assign n2912 = ( ~x4 & x5 ) | ( ~x4 & n1033 ) | ( x5 & n1033 ) ;
  assign n2913 = n2911 & n2912 ;
  assign n2914 = ~x0 & n2913 ;
  assign n2915 = x2 & ~n2914 ;
  assign n2916 = n2910 & ~n2915 ;
  assign n2917 = x3 | n2916 ;
  assign n2918 = ( x1 & ~x2 ) | ( x1 & n754 ) | ( ~x2 & n754 ) ;
  assign n2919 = ( x1 & x2 ) | ( x1 & n1841 ) | ( x2 & n1841 ) ;
  assign n2920 = ~n2918 & n2919 ;
  assign n2921 = ( ~x4 & n171 ) | ( ~x4 & n2920 ) | ( n171 & n2920 ) ;
  assign n2922 = n511 & ~n2921 ;
  assign n2923 = ( n511 & n2920 ) | ( n511 & ~n2922 ) | ( n2920 & ~n2922 ) ;
  assign n2924 = ~x0 & n2923 ;
  assign n2925 = x3 & ~n2924 ;
  assign n2926 = n2917 & ~n2925 ;
  assign n2927 = ( x6 & x8 ) | ( x6 & ~n2926 ) | ( x8 & ~n2926 ) ;
  assign n2928 = x6 & ~n2927 ;
  assign n2929 = ( x8 & ~n2927 ) | ( x8 & n2928 ) | ( ~n2927 & n2928 ) ;
  assign n2930 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n2931 = ( x1 & ~x5 ) | ( x1 & n2930 ) | ( ~x5 & n2930 ) ;
  assign n2932 = ( x0 & x2 ) | ( x0 & n2931 ) | ( x2 & n2931 ) ;
  assign n2933 = n2930 & ~n2932 ;
  assign n2934 = ( n2931 & ~n2932 ) | ( n2931 & n2933 ) | ( ~n2932 & n2933 ) ;
  assign n2935 = ( ~x4 & x7 ) | ( ~x4 & n2934 ) | ( x7 & n2934 ) ;
  assign n2936 = ( x6 & ~x7 ) | ( x6 & n2935 ) | ( ~x7 & n2935 ) ;
  assign n2937 = ( x4 & ~x6 ) | ( x4 & n2935 ) | ( ~x6 & n2935 ) ;
  assign n2938 = n2936 & n2937 ;
  assign n2939 = ( x2 & x6 ) | ( x2 & ~n738 ) | ( x6 & ~n738 ) ;
  assign n2940 = ( ~x2 & x5 ) | ( ~x2 & n2939 ) | ( x5 & n2939 ) ;
  assign n2941 = ( ~x6 & x7 ) | ( ~x6 & n2940 ) | ( x7 & n2940 ) ;
  assign n2942 = n2939 & n2941 ;
  assign n2943 = ( x4 & ~n101 ) | ( x4 & n2942 ) | ( ~n101 & n2942 ) ;
  assign n2944 = n2942 & ~n2943 ;
  assign n2945 = n2938 | n2944 ;
  assign n2946 = x3 | n2945 ;
  assign n2947 = x7 & ~n539 ;
  assign n2948 = ( ~n572 & n1287 ) | ( ~n572 & n2947 ) | ( n1287 & n2947 ) ;
  assign n2949 = x1 & ~n2948 ;
  assign n2950 = ( x2 & ~x4 ) | ( x2 & n551 ) | ( ~x4 & n551 ) ;
  assign n2951 = ( x4 & x6 ) | ( x4 & n551 ) | ( x6 & n551 ) ;
  assign n2952 = ( x2 & x7 ) | ( x2 & ~n2951 ) | ( x7 & ~n2951 ) ;
  assign n2953 = ~n2950 & n2952 ;
  assign n2954 = x1 | n2953 ;
  assign n2955 = ( ~x1 & n2949 ) | ( ~x1 & n2954 ) | ( n2949 & n2954 ) ;
  assign n2956 = x5 | n2955 ;
  assign n2957 = x1 & x6 ;
  assign n2958 = x7 | n57 ;
  assign n2959 = ( ~n566 & n2957 ) | ( ~n566 & n2958 ) | ( n2957 & n2958 ) ;
  assign n2960 = ~x4 & n2959 ;
  assign n2961 = x5 & ~n2960 ;
  assign n2962 = n2956 & ~n2961 ;
  assign n2963 = ~x0 & n2962 ;
  assign n2964 = x3 & ~n2963 ;
  assign n2965 = n2946 & ~n2964 ;
  assign n2966 = n2929 | n2965 ;
  assign n2967 = ( ~n2809 & n2901 ) | ( ~n2809 & n2966 ) | ( n2901 & n2966 ) ;
  assign n2968 = n2809 | n2967 ;
  assign n2969 = ( n106 & n1596 ) | ( n106 & ~n1731 ) | ( n1596 & ~n1731 ) ;
  assign n2970 = ( x1 & ~x3 ) | ( x1 & n1803 ) | ( ~x3 & n1803 ) ;
  assign n2971 = ~x1 & n2970 ;
  assign n2972 = x0 & n2971 ;
  assign n2973 = n1596 & n2972 ;
  assign n2974 = ( n1731 & n2969 ) | ( n1731 & n2973 ) | ( n2969 & n2973 ) ;
  assign n2975 = ~x8 & n60 ;
  assign n2976 = x5 & n2975 ;
  assign n2977 = ( ~x1 & x3 ) | ( ~x1 & x5 ) | ( x3 & x5 ) ;
  assign n2978 = ( x5 & x8 ) | ( x5 & ~n2977 ) | ( x8 & ~n2977 ) ;
  assign n2979 = ( x1 & ~x3 ) | ( x1 & n2978 ) | ( ~x3 & n2978 ) ;
  assign n2980 = n2977 & n2979 ;
  assign n2981 = ( ~n2978 & n2979 ) | ( ~n2978 & n2980 ) | ( n2979 & n2980 ) ;
  assign n2982 = ~x4 & n2981 ;
  assign n2983 = ~x0 & n2982 ;
  assign n2984 = n1536 | n2983 ;
  assign n2985 = ( n1357 & n2983 ) | ( n1357 & n2984 ) | ( n2983 & n2984 ) ;
  assign n2986 = ~x2 & n2985 ;
  assign n2987 = n106 | n2986 ;
  assign n2988 = ( n2976 & n2986 ) | ( n2976 & n2987 ) | ( n2986 & n2987 ) ;
  assign n2989 = ( x0 & x6 ) | ( x0 & ~x8 ) | ( x6 & ~x8 ) ;
  assign n2990 = ( x4 & ~x6 ) | ( x4 & n2989 ) | ( ~x6 & n2989 ) ;
  assign n2991 = ( x0 & ~x8 ) | ( x0 & n2990 ) | ( ~x8 & n2990 ) ;
  assign n2992 = ~n2989 & n2991 ;
  assign n2993 = ( ~n2990 & n2991 ) | ( ~n2990 & n2992 ) | ( n2991 & n2992 ) ;
  assign n2994 = x2 | n2993 ;
  assign n2995 = x4 & n920 ;
  assign n2996 = ~x0 & n2995 ;
  assign n2997 = x2 & ~n2996 ;
  assign n2998 = n2994 & ~n2997 ;
  assign n2999 = x1 | n2998 ;
  assign n3000 = x2 & x8 ;
  assign n3001 = ( x4 & x6 ) | ( x4 & n3000 ) | ( x6 & n3000 ) ;
  assign n3002 = ( x6 & x8 ) | ( x6 & ~n3001 ) | ( x8 & ~n3001 ) ;
  assign n3003 = ( x2 & x4 ) | ( x2 & n3002 ) | ( x4 & n3002 ) ;
  assign n3004 = ~n3001 & n3003 ;
  assign n3005 = ~x0 & n3004 ;
  assign n3006 = x1 & ~n3005 ;
  assign n3007 = n2999 & ~n3006 ;
  assign n3008 = x5 | n3007 ;
  assign n3009 = ( x2 & x4 ) | ( x2 & x6 ) | ( x4 & x6 ) ;
  assign n3010 = ( x4 & x6 ) | ( x4 & ~n3009 ) | ( x6 & ~n3009 ) ;
  assign n3011 = ( x1 & x4 ) | ( x1 & n3010 ) | ( x4 & n3010 ) ;
  assign n3012 = ( n511 & n3009 ) | ( n511 & ~n3011 ) | ( n3009 & ~n3011 ) ;
  assign n3013 = n105 & n452 ;
  assign n3014 = x8 | n3013 ;
  assign n3015 = ( n3012 & n3013 ) | ( n3012 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3016 = ~x0 & n3015 ;
  assign n3017 = x5 & ~n3016 ;
  assign n3018 = n3008 & ~n3017 ;
  assign n3019 = x3 | n3018 ;
  assign n3020 = ( x6 & ~x8 ) | ( x6 & n589 ) | ( ~x8 & n589 ) ;
  assign n3021 = ( x1 & x6 ) | ( x1 & n589 ) | ( x6 & n589 ) ;
  assign n3022 = ( n1461 & n3020 ) | ( n1461 & ~n3021 ) | ( n3020 & ~n3021 ) ;
  assign n3023 = x4 & n3022 ;
  assign n3024 = ( x1 & ~x6 ) | ( x1 & x8 ) | ( ~x6 & x8 ) ;
  assign n3025 = ( ~x5 & x8 ) | ( ~x5 & n3024 ) | ( x8 & n3024 ) ;
  assign n3026 = x8 & ~n3025 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = ( ~x8 & n3026 ) | ( ~x8 & n3027 ) | ( n3026 & n3027 ) ;
  assign n3029 = x4 | n3028 ;
  assign n3030 = ( ~x4 & n3023 ) | ( ~x4 & n3029 ) | ( n3023 & n3029 ) ;
  assign n3031 = x2 & n3030 ;
  assign n3032 = ( x1 & x6 ) | ( x1 & ~n2784 ) | ( x6 & ~n2784 ) ;
  assign n3033 = ( x5 & ~x8 ) | ( x5 & n3032 ) | ( ~x8 & n3032 ) ;
  assign n3034 = n2784 & n3033 ;
  assign n3035 = ( ~n3032 & n3033 ) | ( ~n3032 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = x4 & ~n3035 ;
  assign n3037 = n1159 | n1502 ;
  assign n3038 = ~x1 & n3037 ;
  assign n3039 = x4 | n3038 ;
  assign n3040 = ~n3036 & n3039 ;
  assign n3041 = x2 | n3040 ;
  assign n3042 = ( ~x2 & n3031 ) | ( ~x2 & n3041 ) | ( n3031 & n3041 ) ;
  assign n3043 = ~x0 & n3042 ;
  assign n3044 = x3 & ~n3043 ;
  assign n3045 = n3019 & ~n3044 ;
  assign n3046 = n320 & n729 ;
  assign n3047 = n37 & n3046 ;
  assign n3048 = ( ~x1 & x6 ) | ( ~x1 & n589 ) | ( x6 & n589 ) ;
  assign n3049 = ( x6 & x8 ) | ( x6 & ~n589 ) | ( x8 & ~n589 ) ;
  assign n3050 = ( ~x1 & x5 ) | ( ~x1 & n3049 ) | ( x5 & n3049 ) ;
  assign n3051 = ~n3048 & n3050 ;
  assign n3052 = x3 | n3051 ;
  assign n3053 = x1 | n983 ;
  assign n3054 = x3 & n3053 ;
  assign n3055 = n3052 & ~n3054 ;
  assign n3056 = ( ~x0 & n3047 ) | ( ~x0 & n3055 ) | ( n3047 & n3055 ) ;
  assign n3057 = x2 & ~n3056 ;
  assign n3058 = ( x2 & n3047 ) | ( x2 & ~n3057 ) | ( n3047 & ~n3057 ) ;
  assign n3059 = n243 & n3058 ;
  assign n3060 = n1553 & ~n2735 ;
  assign n3061 = x6 & n118 ;
  assign n3062 = ( x6 & n825 ) | ( x6 & ~n3061 ) | ( n825 & ~n3061 ) ;
  assign n3063 = ( x3 & ~x8 ) | ( x3 & n3062 ) | ( ~x8 & n3062 ) ;
  assign n3064 = ( ~x7 & x8 ) | ( ~x7 & n3063 ) | ( x8 & n3063 ) ;
  assign n3065 = ( ~x3 & x7 ) | ( ~x3 & n3063 ) | ( x7 & n3063 ) ;
  assign n3066 = n3064 | n3065 ;
  assign n3067 = ( x4 & x5 ) | ( x4 & n3066 ) | ( x5 & n3066 ) ;
  assign n3068 = n3060 & n3067 ;
  assign n3069 = ( ~n3060 & n3066 ) | ( ~n3060 & n3068 ) | ( n3066 & n3068 ) ;
  assign n3070 = x2 & ~n3069 ;
  assign n3071 = ( x5 & x6 ) | ( x5 & ~x7 ) | ( x6 & ~x7 ) ;
  assign n3072 = x8 | n3071 ;
  assign n3073 = ~n607 & n3072 ;
  assign n3074 = ( x3 & ~x4 ) | ( x3 & n3073 ) | ( ~x4 & n3073 ) ;
  assign n3075 = ( x5 & n49 ) | ( x5 & n145 ) | ( n49 & n145 ) ;
  assign n3076 = ( ~x5 & x7 ) | ( ~x5 & n3075 ) | ( x7 & n3075 ) ;
  assign n3077 = ( ~x8 & n49 ) | ( ~x8 & n3076 ) | ( n49 & n3076 ) ;
  assign n3078 = ( ~n49 & n3075 ) | ( ~n49 & n3077 ) | ( n3075 & n3077 ) ;
  assign n3079 = ( x3 & x4 ) | ( x3 & ~n3078 ) | ( x4 & ~n3078 ) ;
  assign n3080 = n3074 & ~n3079 ;
  assign n3081 = ( x6 & x8 ) | ( x6 & n357 ) | ( x8 & n357 ) ;
  assign n3082 = ( x5 & x6 ) | ( x5 & ~n3081 ) | ( x6 & ~n3081 ) ;
  assign n3083 = ( x7 & x8 ) | ( x7 & n3082 ) | ( x8 & n3082 ) ;
  assign n3084 = n3081 & ~n3083 ;
  assign n3085 = ( ~x3 & x4 ) | ( ~x3 & n3084 ) | ( x4 & n3084 ) ;
  assign n3086 = ( x7 & x8 ) | ( x7 & n597 ) | ( x8 & n597 ) ;
  assign n3087 = ( x5 & x8 ) | ( x5 & n597 ) | ( x8 & n597 ) ;
  assign n3088 = ( n130 & n3086 ) | ( n130 & ~n3087 ) | ( n3086 & ~n3087 ) ;
  assign n3089 = ( x3 & x4 ) | ( x3 & n3088 ) | ( x4 & n3088 ) ;
  assign n3090 = n3085 & n3089 ;
  assign n3091 = n3080 | n3090 ;
  assign n3092 = ~x2 & n3091 ;
  assign n3093 = n3070 | n3092 ;
  assign n3094 = ( ~x0 & x1 ) | ( ~x0 & n3093 ) | ( x1 & n3093 ) ;
  assign n3095 = n26 & n584 ;
  assign n3096 = x6 | n1644 ;
  assign n3097 = ( x6 & ~x8 ) | ( x6 & n1644 ) | ( ~x8 & n1644 ) ;
  assign n3098 = ( x8 & ~n3096 ) | ( x8 & n3097 ) | ( ~n3096 & n3097 ) ;
  assign n3099 = n3095 | n3098 ;
  assign n3100 = ( ~x7 & n3095 ) | ( ~x7 & n3099 ) | ( n3095 & n3099 ) ;
  assign n3101 = x2 | n3100 ;
  assign n3102 = ~x8 & n218 ;
  assign n3103 = ( x3 & x4 ) | ( x3 & ~n3102 ) | ( x4 & ~n3102 ) ;
  assign n3104 = ( n218 & n3102 ) | ( n218 & ~n3103 ) | ( n3102 & ~n3103 ) ;
  assign n3105 = x6 & n3104 ;
  assign n3106 = x2 & ~n3105 ;
  assign n3107 = n3101 & ~n3106 ;
  assign n3108 = ( x4 & ~x6 ) | ( x4 & n1644 ) | ( ~x6 & n1644 ) ;
  assign n3109 = x4 & ~n3108 ;
  assign n3110 = n3108 | n3109 ;
  assign n3111 = ( ~x4 & n3109 ) | ( ~x4 & n3110 ) | ( n3109 & n3110 ) ;
  assign n3112 = ( ~x2 & x7 ) | ( ~x2 & n3111 ) | ( x7 & n3111 ) ;
  assign n3113 = ( ~n1803 & n3107 ) | ( ~n1803 & n3112 ) | ( n3107 & n3112 ) ;
  assign n3114 = ~x5 & n3113 ;
  assign n3115 = ( x3 & ~x7 ) | ( x3 & n1885 ) | ( ~x7 & n1885 ) ;
  assign n3116 = x2 & ~n1885 ;
  assign n3117 = ( x8 & ~n1885 ) | ( x8 & n3116 ) | ( ~n1885 & n3116 ) ;
  assign n3118 = n3115 & ~n3117 ;
  assign n3119 = x6 | n3118 ;
  assign n3120 = x7 | n1784 ;
  assign n3121 = ( ~x2 & n1784 ) | ( ~x2 & n3120 ) | ( n1784 & n3120 ) ;
  assign n3122 = x3 & ~n3121 ;
  assign n3123 = x6 & ~n3122 ;
  assign n3124 = n3119 & ~n3123 ;
  assign n3125 = x4 & n3124 ;
  assign n3126 = x6 & n261 ;
  assign n3127 = n68 & n3126 ;
  assign n3128 = n3125 | n3127 ;
  assign n3129 = x5 & n3128 ;
  assign n3130 = n3114 | n3129 ;
  assign n3131 = ( x0 & x1 ) | ( x0 & ~n3130 ) | ( x1 & ~n3130 ) ;
  assign n3132 = n3094 & ~n3131 ;
  assign n3133 = ( ~x6 & x7 ) | ( ~x6 & n3009 ) | ( x7 & n3009 ) ;
  assign n3134 = ( x2 & x4 ) | ( x2 & n3133 ) | ( x4 & n3133 ) ;
  assign n3135 = n3009 & ~n3134 ;
  assign n3136 = ( n3133 & ~n3134 ) | ( n3133 & n3135 ) | ( ~n3134 & n3135 ) ;
  assign n3137 = ( x3 & n1484 ) | ( x3 & n3136 ) | ( n1484 & n3136 ) ;
  assign n3138 = n3136 & ~n3137 ;
  assign n3139 = ( x3 & x4 ) | ( x3 & x6 ) | ( x4 & x6 ) ;
  assign n3140 = ( x3 & x8 ) | ( x3 & ~n3139 ) | ( x8 & ~n3139 ) ;
  assign n3141 = ( ~x6 & x8 ) | ( ~x6 & n3139 ) | ( x8 & n3139 ) ;
  assign n3142 = ~n3140 & n3141 ;
  assign n3143 = x2 & ~n3142 ;
  assign n3144 = ~x3 & n1384 ;
  assign n3145 = x2 | n3144 ;
  assign n3146 = ~n3143 & n3145 ;
  assign n3147 = ( ~x1 & x7 ) | ( ~x1 & n3146 ) | ( x7 & n3146 ) ;
  assign n3148 = ~x4 & n10 ;
  assign n3149 = ( x2 & x3 ) | ( x2 & n3148 ) | ( x3 & n3148 ) ;
  assign n3150 = ~x2 & n3149 ;
  assign n3151 = x1 & n3150 ;
  assign n3152 = ( n3146 & ~n3147 ) | ( n3146 & n3151 ) | ( ~n3147 & n3151 ) ;
  assign n3153 = n10 & n99 ;
  assign n3154 = ( x4 & x6 ) | ( x4 & n3153 ) | ( x6 & n3153 ) ;
  assign n3155 = ~x6 & n3154 ;
  assign n3156 = ( ~n3138 & n3152 ) | ( ~n3138 & n3155 ) | ( n3152 & n3155 ) ;
  assign n3157 = x0 & ~n3155 ;
  assign n3158 = ( n3138 & n3156 ) | ( n3138 & ~n3157 ) | ( n3156 & ~n3157 ) ;
  assign n3159 = n3132 | n3158 ;
  assign n3160 = ( n3058 & ~n3059 ) | ( n3058 & n3159 ) | ( ~n3059 & n3159 ) ;
  assign n3161 = n3045 | n3160 ;
  assign n3162 = ( ~n2974 & n2988 ) | ( ~n2974 & n3161 ) | ( n2988 & n3161 ) ;
  assign n3163 = n2974 | n3162 ;
  assign n3164 = ~x5 & n525 ;
  assign n3165 = ( x2 & ~x3 ) | ( x2 & n3164 ) | ( ~x3 & n3164 ) ;
  assign n3166 = ( n525 & n3164 ) | ( n525 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3167 = x1 & n3166 ;
  assign n3168 = ( ~x2 & x4 ) | ( ~x2 & n1398 ) | ( x4 & n1398 ) ;
  assign n3169 = ( x2 & x5 ) | ( x2 & ~n3168 ) | ( x5 & ~n3168 ) ;
  assign n3170 = ( n37 & n1398 ) | ( n37 & ~n3169 ) | ( n1398 & ~n3169 ) ;
  assign n3171 = x1 | n3170 ;
  assign n3172 = ( ~x1 & n3167 ) | ( ~x1 & n3171 ) | ( n3167 & n3171 ) ;
  assign n3173 = x8 & ~n3172 ;
  assign n3174 = x1 | x5 ;
  assign n3175 = ( x3 & x5 ) | ( x3 & ~n3174 ) | ( x5 & ~n3174 ) ;
  assign n3176 = ( x2 & x3 ) | ( x2 & ~n3174 ) | ( x3 & ~n3174 ) ;
  assign n3177 = ( n155 & n3175 ) | ( n155 & ~n3176 ) | ( n3175 & ~n3176 ) ;
  assign n3178 = ~x4 & n3177 ;
  assign n3179 = x8 | n3178 ;
  assign n3180 = ~n3173 & n3179 ;
  assign n3181 = ( x0 & ~n2314 ) | ( x0 & n3180 ) | ( ~n2314 & n3180 ) ;
  assign n3182 = x4 & n2560 ;
  assign n3183 = ( ~x3 & x4 ) | ( ~x3 & n2560 ) | ( x4 & n2560 ) ;
  assign n3184 = ( x3 & ~n3182 ) | ( x3 & n3183 ) | ( ~n3182 & n3183 ) ;
  assign n3185 = x1 | n3184 ;
  assign n3186 = x2 | n3185 ;
  assign n3187 = ( x0 & n2314 ) | ( x0 & n3186 ) | ( n2314 & n3186 ) ;
  assign n3188 = n3181 & ~n3187 ;
  assign n3189 = ( x1 & n754 ) | ( x1 & n842 ) | ( n754 & n842 ) ;
  assign n3190 = ~n754 & n3189 ;
  assign n3191 = ~x3 & n1841 ;
  assign n3192 = ( x1 & x2 ) | ( x1 & n3191 ) | ( x2 & n3191 ) ;
  assign n3193 = ~x1 & n3192 ;
  assign n3194 = n320 & ~n357 ;
  assign n3195 = n26 & n3194 ;
  assign n3196 = ( ~n3190 & n3193 ) | ( ~n3190 & n3195 ) | ( n3193 & n3195 ) ;
  assign n3197 = x0 & ~n3195 ;
  assign n3198 = ( n3190 & n3196 ) | ( n3190 & ~n3197 ) | ( n3196 & ~n3197 ) ;
  assign n3199 = n762 & n3198 ;
  assign n3200 = ( ~n99 & n118 ) | ( ~n99 & n2261 ) | ( n118 & n2261 ) ;
  assign n3201 = n99 & n3200 ;
  assign n3202 = ( x2 & x6 ) | ( x2 & x7 ) | ( x6 & x7 ) ;
  assign n3203 = ( x2 & x8 ) | ( x2 & ~n3202 ) | ( x8 & ~n3202 ) ;
  assign n3204 = ( ~x7 & x8 ) | ( ~x7 & n3202 ) | ( x8 & n3202 ) ;
  assign n3205 = ~n3203 & n3204 ;
  assign n3206 = x1 | n3205 ;
  assign n3207 = x2 & n584 ;
  assign n3208 = x1 & ~n3207 ;
  assign n3209 = n3206 & ~n3208 ;
  assign n3210 = x4 & n3209 ;
  assign n3211 = ( x6 & n21 ) | ( x6 & ~n539 ) | ( n21 & ~n539 ) ;
  assign n3212 = n21 & ~n3211 ;
  assign n3213 = n3210 | n3212 ;
  assign n3214 = ( x1 & n3210 ) | ( x1 & n3213 ) | ( n3210 & n3213 ) ;
  assign n3215 = ~n1387 & n3214 ;
  assign n3216 = x5 & ~n978 ;
  assign n3217 = ( ~x3 & x4 ) | ( ~x3 & n3216 ) | ( x4 & n3216 ) ;
  assign n3218 = ( ~n978 & n3216 ) | ( ~n978 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3219 = x7 & n3218 ;
  assign n3220 = ( x3 & ~x4 ) | ( x3 & n187 ) | ( ~x4 & n187 ) ;
  assign n3221 = ( ~x5 & n26 ) | ( ~x5 & n3220 ) | ( n26 & n3220 ) ;
  assign n3222 = ( x5 & ~n1536 ) | ( x5 & n3221 ) | ( ~n1536 & n3221 ) ;
  assign n3223 = ~x7 & n3222 ;
  assign n3224 = ( x7 & ~n3219 ) | ( x7 & n3223 ) | ( ~n3219 & n3223 ) ;
  assign n3225 = x2 | n3224 ;
  assign n3226 = ~x5 & n145 ;
  assign n3227 = n60 & n3226 ;
  assign n3228 = n26 & n226 ;
  assign n3229 = n3227 | n3228 ;
  assign n3230 = x2 & n3229 ;
  assign n3231 = n3225 & ~n3230 ;
  assign n3232 = ( x1 & ~x6 ) | ( x1 & n3231 ) | ( ~x6 & n3231 ) ;
  assign n3233 = n27 & ~n226 ;
  assign n3234 = ( x3 & x8 ) | ( x3 & n487 ) | ( x8 & n487 ) ;
  assign n3235 = ( x7 & x8 ) | ( x7 & ~n3234 ) | ( x8 & ~n3234 ) ;
  assign n3236 = n487 & n3235 ;
  assign n3237 = ( x3 & ~n3234 ) | ( x3 & n3236 ) | ( ~n3234 & n3236 ) ;
  assign n3238 = ( x4 & x5 ) | ( x4 & n3237 ) | ( x5 & n3237 ) ;
  assign n3239 = ( x3 & ~n21 ) | ( x3 & n201 ) | ( ~n21 & n201 ) ;
  assign n3240 = n21 & n3239 ;
  assign n3241 = ~x5 & n3240 ;
  assign n3242 = ( n3237 & ~n3238 ) | ( n3237 & n3241 ) | ( ~n3238 & n3241 ) ;
  assign n3243 = x2 & ~n36 ;
  assign n3244 = n284 & n3243 ;
  assign n3245 = ( n11 & ~n36 ) | ( n11 & n3243 ) | ( ~n36 & n3243 ) ;
  assign n3246 = ( x3 & n3244 ) | ( x3 & n3245 ) | ( n3244 & n3245 ) ;
  assign n3247 = n3242 | n3246 ;
  assign n3248 = ( n27 & ~n3233 ) | ( n27 & n3247 ) | ( ~n3233 & n3247 ) ;
  assign n3249 = ( x1 & x6 ) | ( x1 & n3248 ) | ( x6 & n3248 ) ;
  assign n3250 = ~n3232 & n3249 ;
  assign n3251 = x1 & ~n222 ;
  assign n3252 = x1 | n370 ;
  assign n3253 = ~n3251 & n3252 ;
  assign n3254 = x4 & ~n3253 ;
  assign n3255 = ( x3 & x5 ) | ( x3 & n234 ) | ( x5 & n234 ) ;
  assign n3256 = n232 & ~n3255 ;
  assign n3257 = ( n234 & ~n3255 ) | ( n234 & n3256 ) | ( ~n3255 & n3256 ) ;
  assign n3258 = ~x1 & n3257 ;
  assign n3259 = x4 | n3258 ;
  assign n3260 = ~n3254 & n3259 ;
  assign n3261 = ( x2 & ~x6 ) | ( x2 & n3260 ) | ( ~x6 & n3260 ) ;
  assign n3262 = ( x4 & ~x8 ) | ( x4 & n558 ) | ( ~x8 & n558 ) ;
  assign n3263 = x4 & ~n3262 ;
  assign n3264 = n3262 | n3263 ;
  assign n3265 = ( ~x4 & n3263 ) | ( ~x4 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = x1 & ~n3265 ;
  assign n3267 = ~x4 & n247 ;
  assign n3268 = x1 | n3267 ;
  assign n3269 = ~n3266 & n3268 ;
  assign n3270 = x3 | n3269 ;
  assign n3271 = ( ~x1 & x4 ) | ( ~x1 & x8 ) | ( x4 & x8 ) ;
  assign n3272 = n2755 & n3271 ;
  assign n3273 = ~x5 & n3272 ;
  assign n3274 = x3 & ~n3273 ;
  assign n3275 = n3270 & ~n3274 ;
  assign n3276 = ( x2 & x6 ) | ( x2 & ~n3275 ) | ( x6 & ~n3275 ) ;
  assign n3277 = n3261 & ~n3276 ;
  assign n3278 = ( ~x0 & n3250 ) | ( ~x0 & n3277 ) | ( n3250 & n3277 ) ;
  assign n3279 = ~n3215 & n3278 ;
  assign n3280 = ( ~x0 & n3215 ) | ( ~x0 & n3279 ) | ( n3215 & n3279 ) ;
  assign n3281 = n3201 | n3280 ;
  assign n3282 = ( n3198 & ~n3199 ) | ( n3198 & n3281 ) | ( ~n3199 & n3281 ) ;
  assign n3283 = ( x1 & ~n66 ) | ( x1 & n1368 ) | ( ~n66 & n1368 ) ;
  assign n3284 = ~x1 & n3283 ;
  assign n3285 = ( ~x3 & x5 ) | ( ~x3 & n1808 ) | ( x5 & n1808 ) ;
  assign n3286 = ( x1 & ~x5 ) | ( x1 & n1808 ) | ( ~x5 & n1808 ) ;
  assign n3287 = ( x3 & ~x6 ) | ( x3 & n3286 ) | ( ~x6 & n3286 ) ;
  assign n3288 = n3285 | n3287 ;
  assign n3289 = ( x2 & n3284 ) | ( x2 & ~n3288 ) | ( n3284 & ~n3288 ) ;
  assign n3290 = x4 & ~n3289 ;
  assign n3291 = ( x4 & n3284 ) | ( x4 & ~n3290 ) | ( n3284 & ~n3290 ) ;
  assign n3292 = ( x0 & n21 ) | ( x0 & n3291 ) | ( n21 & n3291 ) ;
  assign n3293 = ( x5 & x6 ) | ( x5 & n321 ) | ( x6 & n321 ) ;
  assign n3294 = ~x6 & n3293 ;
  assign n3295 = ~n21 & n3294 ;
  assign n3296 = ( n3291 & ~n3292 ) | ( n3291 & n3295 ) | ( ~n3292 & n3295 ) ;
  assign n3297 = ( ~x4 & x7 ) | ( ~x4 & x8 ) | ( x7 & x8 ) ;
  assign n3298 = ( x0 & x8 ) | ( x0 & ~n3297 ) | ( x8 & ~n3297 ) ;
  assign n3299 = ( x4 & ~x7 ) | ( x4 & n3298 ) | ( ~x7 & n3298 ) ;
  assign n3300 = n3297 & n3299 ;
  assign n3301 = ( ~n3298 & n3299 ) | ( ~n3298 & n3300 ) | ( n3299 & n3300 ) ;
  assign n3302 = x1 | n3301 ;
  assign n3303 = x4 & ~n291 ;
  assign n3304 = ( x7 & ~n291 ) | ( x7 & n3303 ) | ( ~n291 & n3303 ) ;
  assign n3305 = ~x0 & n3304 ;
  assign n3306 = x1 & ~n3305 ;
  assign n3307 = n3302 & ~n3306 ;
  assign n3308 = x2 | n3307 ;
  assign n3309 = ( x4 & x7 ) | ( x4 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n3310 = ( ~x1 & x7 ) | ( ~x1 & x8 ) | ( x7 & x8 ) ;
  assign n3311 = n3309 | n3310 ;
  assign n3312 = x0 | n3311 ;
  assign n3313 = x2 & n3312 ;
  assign n3314 = n3308 & ~n3313 ;
  assign n3315 = x3 | n3314 ;
  assign n3316 = ( x4 & x7 ) | ( x4 & ~n1328 ) | ( x7 & ~n1328 ) ;
  assign n3317 = ( x1 & x2 ) | ( x1 & ~n3316 ) | ( x2 & ~n3316 ) ;
  assign n3318 = ~n1328 & n3317 ;
  assign n3319 = ( n3316 & n3317 ) | ( n3316 & n3318 ) | ( n3317 & n3318 ) ;
  assign n3320 = x4 & n145 ;
  assign n3321 = ~n15 & n3320 ;
  assign n3322 = x8 & ~n3321 ;
  assign n3323 = ( n3319 & n3321 ) | ( n3319 & ~n3322 ) | ( n3321 & ~n3322 ) ;
  assign n3324 = ~x0 & n3323 ;
  assign n3325 = x3 & ~n3324 ;
  assign n3326 = n3315 & ~n3325 ;
  assign n3327 = x6 & n3326 ;
  assign n3328 = ~n20 & n60 ;
  assign n3329 = ( x0 & x1 ) | ( x0 & ~x4 ) | ( x1 & ~x4 ) ;
  assign n3330 = x0 & ~n3329 ;
  assign n3331 = ( x1 & ~x8 ) | ( x1 & n3330 ) | ( ~x8 & n3330 ) ;
  assign n3332 = ( ~n3329 & n3330 ) | ( ~n3329 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3333 = ( x3 & x7 ) | ( x3 & n3332 ) | ( x7 & n3332 ) ;
  assign n3334 = ( x4 & n101 ) | ( x4 & n1530 ) | ( n101 & n1530 ) ;
  assign n3335 = ~x4 & n3334 ;
  assign n3336 = x7 & n3335 ;
  assign n3337 = ( ~x3 & n3333 ) | ( ~x3 & n3336 ) | ( n3333 & n3336 ) ;
  assign n3338 = ~x2 & n3337 ;
  assign n3339 = n106 | n3338 ;
  assign n3340 = ( n3328 & n3338 ) | ( n3328 & n3339 ) | ( n3338 & n3339 ) ;
  assign n3341 = x6 | n3340 ;
  assign n3342 = ( ~x6 & n3327 ) | ( ~x6 & n3341 ) | ( n3327 & n3341 ) ;
  assign n3343 = n3296 | n3342 ;
  assign n3344 = ( ~n3188 & n3282 ) | ( ~n3188 & n3343 ) | ( n3282 & n3343 ) ;
  assign n3345 = n3188 | n3344 ;
  assign n3346 = x0 & ~x2 ;
  assign n3347 = ( ~x0 & x2 ) | ( ~x0 & n1687 ) | ( x2 & n1687 ) ;
  assign n3348 = x1 & n1687 ;
  assign n3349 = ( n3346 & n3347 ) | ( n3346 & ~n3348 ) | ( n3347 & ~n3348 ) ;
  assign n3350 = ~x8 & n3349 ;
  assign n3351 = n1199 & n1687 ;
  assign n3352 = n3350 | n3351 ;
  assign n3353 = ( ~x0 & n3350 ) | ( ~x0 & n3352 ) | ( n3350 & n3352 ) ;
  assign n3354 = x3 | n3353 ;
  assign n3355 = ~x8 & n1199 ;
  assign n3356 = ( x1 & ~x2 ) | ( x1 & n3355 ) | ( ~x2 & n3355 ) ;
  assign n3357 = ( n1199 & n3355 ) | ( n1199 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3358 = ~x0 & n3357 ;
  assign n3359 = x3 & ~n3358 ;
  assign n3360 = n3354 & ~n3359 ;
  assign n3361 = n754 & n3360 ;
  assign n3362 = ( x8 & n1437 ) | ( x8 & ~n2184 ) | ( n1437 & ~n2184 ) ;
  assign n3363 = x2 & ~n3362 ;
  assign n3364 = x3 & ~n3024 ;
  assign n3365 = n2863 & ~n3364 ;
  assign n3366 = x2 | n3365 ;
  assign n3367 = ( ~x2 & n3363 ) | ( ~x2 & n3366 ) | ( n3363 & n3366 ) ;
  assign n3368 = x0 | n3367 ;
  assign n3369 = x1 | n66 ;
  assign n3370 = x0 & n3369 ;
  assign n3371 = n3368 & ~n3370 ;
  assign n3372 = ( x5 & x7 ) | ( x5 & n3371 ) | ( x7 & n3371 ) ;
  assign n3373 = ( x4 & ~x5 ) | ( x4 & n3372 ) | ( ~x5 & n3372 ) ;
  assign n3374 = ( x4 & x7 ) | ( x4 & ~n3372 ) | ( x7 & ~n3372 ) ;
  assign n3375 = n3373 & ~n3374 ;
  assign n3376 = ~x6 & n145 ;
  assign n3377 = n67 & n3376 ;
  assign n3378 = n99 & ~n3377 ;
  assign n3379 = ( x1 & x6 ) | ( x1 & n171 ) | ( x6 & n171 ) ;
  assign n3380 = ( x6 & x7 ) | ( x6 & ~n3379 ) | ( x7 & ~n3379 ) ;
  assign n3381 = ( x1 & ~x5 ) | ( x1 & n3380 ) | ( ~x5 & n3380 ) ;
  assign n3382 = ~n3379 & n3381 ;
  assign n3383 = x3 | n3382 ;
  assign n3384 = x1 & n552 ;
  assign n3385 = x3 & ~n3384 ;
  assign n3386 = n3383 & ~n3385 ;
  assign n3387 = x2 & n3386 ;
  assign n3388 = ( x3 & x6 ) | ( x3 & n171 ) | ( x6 & n171 ) ;
  assign n3389 = ( x5 & ~x6 ) | ( x5 & n171 ) | ( ~x6 & n171 ) ;
  assign n3390 = ( x3 & x7 ) | ( x3 & ~n3389 ) | ( x7 & ~n3389 ) ;
  assign n3391 = ~n3388 & n3390 ;
  assign n3392 = x1 | n3391 ;
  assign n3393 = ~x3 & n811 ;
  assign n3394 = x1 & ~n3393 ;
  assign n3395 = n3392 & ~n3394 ;
  assign n3396 = ( x1 & ~x3 ) | ( x1 & n572 ) | ( ~x3 & n572 ) ;
  assign n3397 = ( x3 & ~x6 ) | ( x3 & n572 ) | ( ~x6 & n572 ) ;
  assign n3398 = ( x1 & x7 ) | ( x1 & ~n3397 ) | ( x7 & ~n3397 ) ;
  assign n3399 = ~n3396 & n3398 ;
  assign n3400 = n3395 | n3399 ;
  assign n3401 = ~x2 & n3400 ;
  assign n3402 = n3387 | n3401 ;
  assign n3403 = ~x4 & n3402 ;
  assign n3404 = ~x7 & n1961 ;
  assign n3405 = ( x1 & x2 ) | ( x1 & ~n1961 ) | ( x2 & ~n1961 ) ;
  assign n3406 = ( x7 & n105 ) | ( x7 & ~n3405 ) | ( n105 & ~n3405 ) ;
  assign n3407 = ( x7 & n3404 ) | ( x7 & ~n3406 ) | ( n3404 & ~n3406 ) ;
  assign n3408 = ( x3 & x6 ) | ( x3 & n3407 ) | ( x6 & n3407 ) ;
  assign n3409 = ( x5 & ~n105 ) | ( x5 & n1706 ) | ( ~n105 & n1706 ) ;
  assign n3410 = n105 & n3409 ;
  assign n3411 = ~x6 & n3410 ;
  assign n3412 = ( n3407 & ~n3408 ) | ( n3407 & n3411 ) | ( ~n3408 & n3411 ) ;
  assign n3413 = ( x1 & ~x2 ) | ( x1 & x7 ) | ( ~x2 & x7 ) ;
  assign n3414 = ( x3 & ~x7 ) | ( x3 & n3413 ) | ( ~x7 & n3413 ) ;
  assign n3415 = ( x1 & ~x2 ) | ( x1 & n3414 ) | ( ~x2 & n3414 ) ;
  assign n3416 = ~n3413 & n3415 ;
  assign n3417 = ( ~n3414 & n3415 ) | ( ~n3414 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3418 = ( x5 & x6 ) | ( x5 & ~n3417 ) | ( x6 & ~n3417 ) ;
  assign n3419 = ( x2 & ~x3 ) | ( x2 & x5 ) | ( ~x3 & x5 ) ;
  assign n3420 = ( ~x5 & x7 ) | ( ~x5 & n3419 ) | ( x7 & n3419 ) ;
  assign n3421 = ( x2 & ~x3 ) | ( x2 & n3420 ) | ( ~x3 & n3420 ) ;
  assign n3422 = ~n3419 & n3421 ;
  assign n3423 = ( ~n3420 & n3421 ) | ( ~n3420 & n3422 ) | ( n3421 & n3422 ) ;
  assign n3424 = x6 & n3423 ;
  assign n3425 = ( n3417 & n3418 ) | ( n3417 & n3424 ) | ( n3418 & n3424 ) ;
  assign n3426 = n3412 | n3425 ;
  assign n3427 = x4 & n3426 ;
  assign n3428 = n3403 | n3427 ;
  assign n3429 = ( x0 & ~x8 ) | ( x0 & n3428 ) | ( ~x8 & n3428 ) ;
  assign n3430 = n15 | n587 ;
  assign n3431 = ( n10 & n95 ) | ( n10 & n3430 ) | ( n95 & n3430 ) ;
  assign n3432 = n10 & ~n3431 ;
  assign n3433 = ~x0 & n3432 ;
  assign n3434 = ( n3428 & ~n3429 ) | ( n3428 & n3433 ) | ( ~n3429 & n3433 ) ;
  assign n3435 = ( x4 & ~n105 ) | ( x4 & n1420 ) | ( ~n105 & n1420 ) ;
  assign n3436 = n105 & n3435 ;
  assign n3437 = ~x8 & n3436 ;
  assign n3438 = ( x1 & x2 ) | ( x1 & ~x6 ) | ( x2 & ~x6 ) ;
  assign n3439 = ( ~x2 & x6 ) | ( ~x2 & n3438 ) | ( x6 & n3438 ) ;
  assign n3440 = ( x2 & x4 ) | ( x2 & ~n3439 ) | ( x4 & ~n3439 ) ;
  assign n3441 = ( n354 & n3438 ) | ( n354 & ~n3440 ) | ( n3438 & ~n3440 ) ;
  assign n3442 = ( x3 & x8 ) | ( x3 & n3441 ) | ( x8 & n3441 ) ;
  assign n3443 = ( n3437 & n3441 ) | ( n3437 & ~n3442 ) | ( n3441 & ~n3442 ) ;
  assign n3444 = ~x5 & n3443 ;
  assign n3445 = x4 & n1437 ;
  assign n3446 = ( ~x1 & x4 ) | ( ~x1 & n1420 ) | ( x4 & n1420 ) ;
  assign n3447 = x1 & ~n1420 ;
  assign n3448 = ( ~n3445 & n3446 ) | ( ~n3445 & n3447 ) | ( n3446 & n3447 ) ;
  assign n3449 = ( x2 & x8 ) | ( x2 & ~n3448 ) | ( x8 & ~n3448 ) ;
  assign n3450 = ( ~n3437 & n3448 ) | ( ~n3437 & n3449 ) | ( n3448 & n3449 ) ;
  assign n3451 = ( n312 & n729 ) | ( n312 & ~n2347 ) | ( n729 & ~n2347 ) ;
  assign n3452 = ( x1 & x4 ) | ( x1 & ~n3451 ) | ( x4 & ~n3451 ) ;
  assign n3453 = ( x3 & ~x4 ) | ( x3 & n3452 ) | ( ~x4 & n3452 ) ;
  assign n3454 = ( x1 & x3 ) | ( x1 & ~n3452 ) | ( x3 & ~n3452 ) ;
  assign n3455 = n3453 & ~n3454 ;
  assign n3456 = n3450 & ~n3455 ;
  assign n3457 = x5 & ~n3456 ;
  assign n3458 = n3444 | n3457 ;
  assign n3459 = x1 | x6 ;
  assign n3460 = ( n67 & n576 ) | ( n67 & n3459 ) | ( n576 & n3459 ) ;
  assign n3461 = ( ~x4 & n67 ) | ( ~x4 & n3460 ) | ( n67 & n3460 ) ;
  assign n3462 = ~x4 & n1502 ;
  assign n3463 = x1 & n3462 ;
  assign n3464 = x8 | n3463 ;
  assign n3465 = ( n3461 & n3463 ) | ( n3461 & n3464 ) | ( n3463 & n3464 ) ;
  assign n3466 = ( x2 & x3 ) | ( x2 & n3465 ) | ( x3 & n3465 ) ;
  assign n3467 = ( ~n36 & n3458 ) | ( ~n36 & n3466 ) | ( n3458 & n3466 ) ;
  assign n3468 = ( x1 & x2 ) | ( x1 & x6 ) | ( x2 & x6 ) ;
  assign n3469 = ( x1 & x3 ) | ( x1 & ~n3468 ) | ( x3 & ~n3468 ) ;
  assign n3470 = ( ~x2 & x3 ) | ( ~x2 & n3468 ) | ( x3 & n3468 ) ;
  assign n3471 = ~n3469 & n3470 ;
  assign n3472 = x0 | n3471 ;
  assign n3473 = x3 | n1287 ;
  assign n3474 = x1 | n3473 ;
  assign n3475 = x0 & n3474 ;
  assign n3476 = n3472 & ~n3475 ;
  assign n3477 = ( x4 & x8 ) | ( x4 & n3476 ) | ( x8 & n3476 ) ;
  assign n3478 = ( x5 & ~x8 ) | ( x5 & n3477 ) | ( ~x8 & n3477 ) ;
  assign n3479 = ( x4 & x5 ) | ( x4 & ~n3477 ) | ( x5 & ~n3477 ) ;
  assign n3480 = n3478 & ~n3479 ;
  assign n3481 = x0 & ~n3480 ;
  assign n3482 = ( n3467 & n3480 ) | ( n3467 & ~n3481 ) | ( n3480 & ~n3481 ) ;
  assign n3483 = n3434 | n3482 ;
  assign n3484 = ( n99 & ~n3378 ) | ( n99 & n3483 ) | ( ~n3378 & n3483 ) ;
  assign n3485 = n3375 | n3484 ;
  assign n3486 = ( n3360 & ~n3361 ) | ( n3360 & n3485 ) | ( ~n3361 & n3485 ) ;
  assign y0 = n35 ;
  assign y1 = n110 ;
  assign y2 = n212 ;
  assign y3 = n329 ;
  assign y4 = n518 ;
  assign y5 = n737 ;
  assign y6 = n919 ;
  assign y7 = n1094 ;
  assign y8 = n1286 ;
  assign y9 = n1479 ;
  assign y10 = n1665 ;
  assign y11 = n1855 ;
  assign y12 = n2045 ;
  assign y13 = n2211 ;
  assign y14 = n2409 ;
  assign y15 = n2578 ;
  assign y16 = n2774 ;
  assign y17 = n2968 ;
  assign y18 = n3163 ;
  assign y19 = n3345 ;
  assign y20 = n3486 ;
endmodule
